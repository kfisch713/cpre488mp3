XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��L�JH��0����@8�O��'A3���(��ຽ#^�/�ӎS�&|�榙=��z���k5����Eק���%�g�%LsS�B�A�}�na��j��_�v�K��[a�$$6��).�9�J�2�١)���@di⠺��������	˿��@=[C��8s·�� �8�c0�G&�k��5�ٝ�|�z?x�qx�J�t���7�_���7����;����)N%��K ���c���=��8�x��%���*�Q��R���I�F�6�K�#%C,��f�����ɜMв�� �ڹ<�D��Y�ϓ�@3g���ۯl"p�h�[Q�oC{�"$4W��v�ʄ
r������|KMaXs\]�����oI������T	�o�߁ç|�:wx���-��eiU�R¦���
F�I��S�\�+�Y��X�8���B�1f��� ���5���:��Ϸ]���r���Ud֑�1���~F��7RQ+��2�~��"M4?ۭ��B���hNg�e�W��[o�E��	v�tR=�y�A"��в�r:��0�zR���[��8ӑ��~W��d0R]}<i"�,��{Fi��K���SRPw�X_ "WaY�m���S�u�fɪ���/�X����B�!+D@����Z"��,M��.E�t����mO,�d�� ��/* }�)������ڪ̿հ��wF`/�(���BA�`���x��!�����������2� ��Ԧ(W���X��`q\_�XlxVHYEB    1448     800�Or��d�f�!�0����X�@q��ׁ��H��0d�T�6�lڙ�}��������}��L��&ZU�}��sۉT3_t�KQ��+Q/�8�� �Ć��@8��0��*��|��K9�U{���w�a�Dh��ƣ8^$��ߺ�ø�o2a�<L{XWY[�+%7��-���}��Q�y�֣�؊��ӛӌFU�0��v`?-N��i>�B�mK�΄sM}�<X������xX��R��)<�{�hz�'�ˢ	�+���k���ۣ����{D�-oi�	y	�O�?e���~�2O�߫���K�9�n�O���'<"រ��70��r�"O�M���#R��mn�Rܤ�,%�+L(��<(�ӄs ���6�_ �a�9�,�a/k��26�7�P��T�xJ{�L9�ӟ�=�[�F���ia������c;���Ç��3m[\pHՏ�JD���ю���ڡ Q�rOp#���˟��1�8_N�i�?�̃@�Y��&��a�H������\A>.8緎&���~�8��0�0�b����N�5��ͬ]ҵP[2�;�-F�%p!E�d����/ ��{Ǯٚ��^G��%�{v� -.�8H�Śg{qO���+W���+�|����(a����WeR�8�H��\\��bPF�h��Q*�+P�A��4��Յ�BR�I�M���'D�4��6M�n�ǈ?j9�8O| ��i�m��)I��D��M����`1��G-_ X��(-t+r�������Q�"�z�l56 ���Y��>b���a���I���e��׊�t���!��j��Zؽ�����ۃv����L���������ڹ�Ƭ���n�O�5�p����&�wv�N(Y��k�b1_��G��1��n9M�2�*�C��ʗ6f;��E�H�vAp>���[�6��i%�m��M�ݫ�ؚ�}��Z=3���Kf�G��B�����e�SN���g-q�{Xڤ],B;qgT��a�����:x�QSV=JF= %q�<��!��
ӟu�=n��χ�m����\�Y=�XdxA#�5����E�v�oޝ�L'�zc����[���f8n�qY
�\�9�cƚ�&#�3�?�OQπ�!���ɹ
0��bO2i�����g�d�_�̕���JP)���c���Oڮ��@�#~��I�&�Ӕ�n���3)�������Ⱥ^�٬��ă�9���P��0�1�Q���r��鷤�q֖�{-��qf'�w1XD+*����j���{4�k%8\��.��蛯����J��|�M�r%Ď���MNz�Ǝ���G}>�S�T���u��/$�¯^��こ�N�V~d�5T�國�,Q��Uؿ.j��rR�=���E���{^�g�Z��m�|�q�:Eh�ҖǨb��>(T��m����o}%�ˊ��Gt0!��9��W.�eI�w�Y��e�@�O��Q�B�q�*q��{�rQ
2��f�DE�MIřk�P`#�*�>�>�U:������T�p9���LQs���*��.����f�:̮ƖRkH����a�zB���aό�*��\?r{�K������fO�_��I�9�Y�DLt��U	y�tx4AG�5|rJ�Y�?Mz
4�ƥ-����,r���W�B�`s����ע�.�j�{s�h�b��߱'�D+�i�������L�p!	3������ѱz��v}E����<��d�W�.7p�kk������v,n�"e(j^�5�Q�z��IjB�|̰~a�s����uΤܢ��ƹ�����	0h�,��\���E�]�.�m�{$[2�g�M������9|�_�j�痶�i`�lXv,�Sc�E �ʵ?�_kx#�xn���:����8�Z��ȖMRuP��<�}�o
f*q��0�?=3SPl�|؀-m%M�_���%�)tv�k"�]��<�2�q9�E�*tq]q��!K���b'wZ���nB��%�Aή�7��C��gՐ�֌ +n�r��#/`,����/� �7�6���F�