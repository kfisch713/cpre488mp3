XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���P+1Cz�R��,���h�W&�*�Z%7�e����}��H:��2ȮM���qH<�G��X���LH7�g��m̼�S�{�Kƶ����;��D���GL%~g^.��:Q�FF/|\��X7NaV��!��t�1��b&y���Ns�g�g}z"L�k�W�c�#�ݗ�h��]�P}����l�q�q����ڿ9��M�~k���ϯ��݊��Sx���9���|�_-u�?��i����^�Cr�s��'T�'�H�*��6zPA�!0������V.�i��~󔅶ы�~��=q��.��u�#����4�//u(�Y�<R�Dv�۱yO�ނ� ~�����u,&c=�kg����F���j�#
��+QH��XquwX@��뢀�LC<��P���Qăֶ�.;�ua,��q�O[x\�ihw�d�|Y�
u_{��o'��I{JxP(���6����Il%������	�q��������^��:�6�\�%I��o$��9UD�/��p=��;���'hW�4ޙ��@���[!�˸ۜ2R
���1ӄ��G�WEe<��F�EO	ⶄG��@K9�X?ge(���#.]�`���h�����J�r[_�E���j���������oI��E# �(��߄�"��x`K�AR�jB�����2�Ɣ�Ł���x��XgI�jy��7aK�.�	4�5�ңР�ZZ`��&^>��d3��=��E���ךiO�Ø��>C"}���\@��P/��eU7������#
3㪤OXlxVHYEB    1853     810���H�6(���ജp���e��%�N����Cw�i(���A�4���RR��K�w�y8\��\6�5w^d�>����ߞԃ���l�u>3�)ʠ'����g�˪#�az���I�P\��BX+���9P��v(
I�?�BPr^�7���*!P����B]X�kI�Gl�刢T�.��X�6�B�
:�DnE��)Sl��=�I����~Vo�CM�������C(�!�k#����F7�g�rr:��$���]��X wvdpF7T���(J����k^X�z�w �1��O�2�;����p�St �&}��͙^zL��v>zP��!Գ�3������X����b����4�k%��z�ǣ��}_��P�@���VC9��+B�a�-� �u��Z �"A6� f�pG��o˜PJS�}P���n�Cߴ���vˠOҖ��+ˈ�Z�)��Ř�`���D���?E��F��(� 	���`��Q[Ѯ�8Qi4���;���Y�T��!H��p=ED�	����Uu3�^�;�uI?5�x륂�sǎ�J6��VD/$���=Ru�%�~b�j𩎮��e�uP-�s�p������:���v�pzoF�MK-\���J��/����l���o!���DR�$**�X�|w��9�]��-�J�M��!͕Ƞ#"�fC`b��f$�����6��a`��μ����v�� ~�m�@����G�Q`���� 0w��M=��
�J~-)	���C	ksG��VLP����g�Oj�����`
����7�>�,#]��t��Fð���]G��.5;��)����|�������X��.��9[���L�>��b��#�@�����I)Qi�~�u&��`�6b�[�O})<�A���x^���˂�;�l�!l�+/�"�CF��
C����j���̨Wc�<H��Y�_0�"#uae�.�T��w( �
ڪ���C�fc%q�bV�t��W��R�j���W���1��{�_y�'����w�v'π���,��=���d6�䑟B��T	E�|e�ڪ><}��1Ň�/���s|��lJ�9�U�]W�!�,���������޴�_5Rx��Uc!
�&�ۖ[āG�"���>V���Z�g9=B^J��y����a����?؟��Gf\��
�_��RH�-�gN�*j[A>/�}:kh1��E�I����xȒe��P"���n�CA���*6]{��X����	\�����@��~*T�M�[���	�<���ѝV'��!
Ѓ@�T�k��r���[[�݌���"�	�+<�ݲ�R�d�j�!!cX�뒯d�AۙP(�7m ��e�u��o�����`�ٺE�+�3�_e�3�`�N��o�2����2��Y�N"�	���H��4�'�Sa~� ���o���ze�0������ܞ菔mՓt�@�m���5�;xg���`?S��(wH$J�����(��?�m�h���^��I�[fBFP�Dۣ�k�ۺ�L��&f�E�SW�\��MF$u5�3�'Y�_��	T{>3衷��pr@�s�q3!��a�^�f;嶘�Л�7d�i���!����J�ǸmuB/Ǹ�I��6cX��7ř�N{�\j�8��AX�\-�FYӜ{fڧP��b��?���2���)��f{�����v��!����!puC"m�'��KP�&C �q����O�jl"��Y�_p�Y_�ߖq�i�G}��מb�����JY1Π{S �m��������G|�����U���	�(���tJW(�=-h����4>DP �If#x�Щ�JMb��3"�@"�^�#�?Z�%�Zg11#��D�?�ثq�=��gǣ��`r��}���F9�W�f�=V��!�Z:�����iE�Y[Q�E�����1m'#��b�B�\�����Y�KZ�k5-ƕ6��-��p|Q�y���>"�w\/Pd�/z5y�:���V7�BO?�C�Q�\��Ϩ�/���Y��ȂJ���B�-�h�޹K��߁� �l�*�sg,r�<