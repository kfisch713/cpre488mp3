XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ѧ�H��- ��R�54W����D��s<���픶�چ�����I��YK���N��-5M��Km�%�K����ۑ���ڐ�2�v/��������]Ψ���Q��4���2Q�F._֕$�D��d�N�d��y�ݶ��_9��p�f�Jq[�����u�1'(p��b6Y���T�� 	W���
�Fj���t S"��F�c"H ��:B�m%2C�4�>�F���m�a�gj|��r�W���p|�ݩ��7���
��|�kŲ�g)�6]Р��ui��4Uàa��M���YE+]��=����^�x�@$ }1�� �lhh��W��hɵ�A!��ė��u�4A��
�f--�ÌF�A��H�v�{Ԁ1Q�$h� � 4m��[v��������c ���]PxWL&�3�B���ej��l?%s�'0�������dM-��(��e�-�!~��O��~W�[�|��ſ�C��襸G�}h=U_r��7�-���.P�f���W�jY�wk))�/���~���M8q簨�O���/�w�N���3���޶��Ql�W�T�@�!�y��~#nf���� �����<.S�Ǆ郷�����0^m6�� ���5]�~�Ӄ�2N���{��4܎9�ȳAMko�5��__Ŷv �Ϊ�����ykkN��?g�6ߵ��>�7���̄���z��dkpO��'vn�~�&}��H�.EÛ9��*���9hV�1|<:��#�9EU�
;�=k�����XlxVHYEB    3da6     fb0r��?/+�i� 1h��L���I�#������j#��E6ܬ��i;���bK�[q[iIGG�֖%��fWQp�M�|�p�)a�j���!' �uկrK:2��Fe���Ѵ�Q,"�z�I�>D��A�CC���"K?�(�7���<�%��Ve�@��%)`�<��7��ܒ���:��呥T�I$�JZ.����R���E�`�&�FR�E>e6OO�Uf��*B"��%-��v��㠂RR�,r�w|0�/�EO,}C��W���4�?M�v6[���W��n��Ep��H��`q�-"x^	aJCE���v�)a��w+v$i����s�+R`��2�Wl�=����(:l�]l;l����0.�'�E�!E{��U�9ċ��TL�����<ױ7��DYs�Ojz���@��^��P䪵�|} :�$'�f�}w��v�s���T���ek��G���0��\�*�lSyR�b@��(%�����-�02V!ZC:�E������w�&ݼ�*8��/�mhC��'�0���8,Jk�Us�~�H;�a��pZjzɈv.�Il5�h�f+H�O��=���Sl�1hv}V\�[N09�䃟a4�@J��C/��B��zU���ԫ�#������	=�az�b���ZK����W��6�|�=��Ά�,��C�.�?z�\���hx�Q�b� �g��%������ ����&Q*��L��ډ�㋔&�Yܶ��  ��7t�GZdO�P���u��C9��T�a�FV[[��zi},/>P�w+z�Ԓ��6R��؜��<8�ڬMU�лGua�0U9�v��e4��V�M�>��m���az��F��V���x��DW��'�q�R~��č����H�u�Үq�����އ�B�"`DDˆ=�oG��̄VR¡S2��Y8�6қF�wP�����f�UM�B�4Z�Sٶ�3�ud�,����xI^hM����.x8��t����p�$�CJU�F���������K�N쀟�[6��." 'P8�{�ʁ��j6�bP��U6K~(�v^)��W�|��L:u���h��0�ѕO���i��8�ƪ���~s�U��^uL��+I�!D�T^����*ޅ�#Q��-�h�p�P�w����SZt�3����tKvr�͉��'����&��δ|$s�m~jnT7λ(W@\a�o0Bɗ/�	l['�D�-��"YY�w,��Z�XŮ4� �*����e���@����v��迁FP�(lɊi/��Q-|�2��^WPL ���LF�ET=Yp��g��g%�e|�Y9mWce�g���z�BpO6�]e/�ʆ���u��\׹`�_�y���^|'��������1Z�r�,��	�����a�qOۅ"�����*�x=#ђ(��1��.�,�x�
�T���9�(詔3ZW�%��ۇt�S�<���C+�N����_���q92� w�rG����N���4����H��c�>�f�����3�����<�f�Vщpm{�U�޻t<;�f~w�dK���7�Q��s�S����d7�^կ��R�+�[��8w3&n��35g�s�u�hB��%#m"6l)��s]�O����P-ϕPVS�~�`Sy�k᪉�+ql'Q�b��Y{�<g���3M�+���`+�8��Y�G���NJSײ��n� l1U5��Z!�܆�Z]nL��k�՚��A^�7�Sj^y���M.=�>Z|��eN&�RÏV���a�����h#����o�6`�(���#XjO\�D+;ưu\�Į���d7 !L'0d��~�ʮ�Z� VԦ]؏{5��T繓dYY��I��ܲ�AO���4
�ߙ�4?e����⻱@����㣁�,{'>�p}����N�'�����呹�H���1��N��
�7H�P74s���O���t6����/o���"�ж�ET�ep�w��_b@ܧ�d�*�A|���W�!$�.T��f�Y��������&;z��7�����o�u���B�B�{�G��lKO�[Pp�^	�7�<N�$�ی�/l��pC����
[�'��:ۅ�NMق
�o�A�#��#�'����dV��T��4�I�L7'�dX��_s���T�3c>2`Hs	k�c�v�4�I��惤{�y�Rw:����C�Y�U�����X��U
E��?Ѻk�����G�s>����BJ�����C�
ii���U�k�?��?Fދ�i�֮�tW/TK�5�t����\QeP�:�����j�\��x�m�R3��I;D4�c�o8�"���ϛU�4��0L"{�P#+?bk	��s�q-)��/��u5��}2�Qk�(a�
1a>���խ�,���p�OT��D胣 ���\���~��C��r���((��S@M���l�ނ�c]��ڒ�GM��� �����]�|L� @VQ���v�hL�m��[S,"	�?�Ԯ��߹RΉԢW-'�!%NZHı(gh=ã����l�!ɵqj��G;�C��7��J�U;Þj��������j<�RP����9����y֔z]f)��%�&��G�]������
��V>3�O��~68��|��%4] �{�M�Fe�)!��m>غ��b��Y'��/�S(Ws�dsck��y4�tۂ�*��iM�I���kK�3�(�x�̃��O�����W��`aNm�_��֒?���1���w�X��u�:����ݲz���@x3h�ƛQ��U� �fل��Ir̡�Ɠ]�&����ҝv��u˦�z�T�vn��I|�/,뮥���<�UPߗ^N6cQ����ϔJ2S�#X�6�����l����6{���+ix�r�є��۱8|��L��-�)��0[!i9Es��mA��/� ;VS��!��2��%^D{�!P��=ǣ��$$pC���V���߻��5�Z���3�B���E�U�ڐ�1�J��˓H#���谁�g�b��a�Q��|�=�v�V�$�!�?�A(5P�F3�H��
���F`�q�_eڥJ���:J�v��zkͻ�8�~�&�a:�����>��,)`�Eb�$���k�I�+��`��Q,���}��<s�X�Q��Qz����u;2�rBC�{r�3�#���:�(%ܰ7��y�5 DP�r����>��^Sm,��� ZI��ʖ�ˑ���Qz�V�Զ�(}5
�� �YY��y�f�"��|I<}Nm�e=�d�J�_KS�C��n@���-�ⷣވa�DSi[Ֆ�ι�@���a�'ME�%\���@WYt0��NN��-������EJ��xR]e����8�^���G�SoY�%(��'IB�4jIԍ��Gڸ`�20�1۾��޸sw�)�E%�0` ����-x���f�"��ʴPOr�3rϡ;5� �w�nC�tDR.ض�ܲ6)���ۃQץN�4#&ط���!6)}:* �PA0�F5J�j$30��{,�pe����'��tg��c���6*_�L�bWD;�X����n$�/Yۏ��/ۨ�k~@�$��f�	�]�;�l��򶑸Q�<~to�)�fhW�\��`"�z(��0���]�=ٻIg��y]�N���5JT��}��1������s
�)�L ^WGY�"����S�	�M���R��?hP�F:���AX�H��bp�Q9h�E?�n�@R�h��`��������Eb*=�;�XYAMpF��\IJ�.�.O㰆���sυ�R��������d���k�p6��~�H!6��g�f��@'&k�{�=��~��Y/	)2�G0IJ0)�Nz��G&�~_�KB���`�v�g��U��ҋ�鹒�⽣�/���C �2&�!#�~��S&���1z�<�AX��PP|�����o����Y�>�l-ޟ]�}ҥ�f�1Y\4D*�Z�c�I