XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��j\�M������hhhfazQ[�����n��b֊�� �)��{�Rc��һ1Gl�<�jX�k.�0���kF��i�8<�F�ng����9ē��
Bqb�%�u�hēd���O��O�2�U��s����sSg�h���M"B�R��-��֞tl�QTTr�&�Uck�^��ʠh�1�OsL�ێ};3�x�Fld��K�%�{Dyzr= �X����ƛ����:\< ����r����8�H���9WK[3DDAH�g�3�B�+;jKzF�c�fSw7�E��yXDN]3��Jf����9g�ؼ��G�k��u�*�`��j������p5��E2�:T�?T�J�<�c��8�(Q*���T���@�]�`A�X�����p� ��|�0��Fϰ=gt��zofv����9�U�Ƃ36ﾣ��;�G�"\��I
!_:=ٴe�����`d��p��gD�ė�?)����	s�p;J�'�� 4=i����6�3����%q���$�G�H���4'��'��Nt�e���t���s���&,���-�>`�@V���T��R�E�%E�t�Ȭ�H��gS}"Oi!�zÕ�P��g.6�����6� ���1a�K�b��ܐ9XƼ�NRt���#_�������۹]C���&�$eM@ ;rL���s8�JZ	�����N퐼�vݽEx{�<]��'�4��r3%�
���'ʾ�XS�Q%�W��w����Ar��Y@��NhZ���2����]
�?����XlxVHYEB    1853     810E���AK�w� ��a��4D�)(�.a�](�
�o]�����$����)ӔP*!ꏓ� {��8�JH��@��KG�,�Ly����w���60���-�5�9�!�v�hc���L`��"N�q��S��逥.�x"�E4��*�DRe�wVG3�J[0�o4�`�A������5LLͥ�>St9N�7��,+���w�W�d�$�l���~p^y(W/����Ս�o.������xX����A +�ؕFe`\�W�%I�Ȇ5x������W;vF-z�����A�ֈ"��J�9Đ߃��0ɦJ[`[��GZn?)?�VdA=c�ngp�4�v�Y��`/�^�g�0Ap����x��zx;t���<��YG���U-�� W���q텇2v��laP�G�
&���Մ��'Tq���!�H�1�z�s+K�5��$�C������/e�Е���<6F%���m����j��iRk��0�������)X�y��,S�c��G��%�@������s�Z�*��1q�Ji�$ ��0�y�9r�s�\� ���y����@���z�P��@Fv�ޏi]5A>�K��0�Wڔ�!T��qJf�B�<��XV��iډ�T�;�Y�\3<!����nZ �\�xjI&X��+qy9&�YK��]�a`��T�'q��oM�	��N)j	Y�C�ߏ!���P�.A@vT�css��'�s�	��\���Yux�n����X��u��V��Ԯ���'�@�=0�y��-�ه�{֤bL�IV�9��&�:�
��T���',��3�sɕN��u��d�Cɛu5&Kb�IWE׬�u�Բ��/��1��u�e�jЪ����O�FCZ/��ܾ�`�<�is�g�M��'��ܮ�M4x�֤�ƫ�8�S\��c���*���$ ؿXڻ� C
�.�ެ;�;�ԉ�M���ҷ	u>�[-b�k�RS��M��_a:h#Qw�j����uYz-[��^nk�j��렻�;�!�^����	!����N��u����ÉsgO�v~^ ��/G�.����D<N5܈oѝ�����./�=�-u�AT��&�
͖���պE�VR�����&1ϙ#N>t��.�gHH����Dz}��3���eL�}R����{���xO�o��]�oe?U&K��v�`[��~�V&8�d����a9	��fB������[��)0w�pVA?N$b@ha+p<��'��NcS�(/ ���P�������ʪ�Z]�P���$�a^Д�n��֙�;�1~���r��o��&a�Wpt�x���E銉|`*y�M��M˲�e�\�"}��r[�}�h|bF�\6T(* *�
���������� �V�XB�K�tu���x�����$�-�G��1�G�<��*��9�l���Qx��٫!���d䧭�yBu�z��̍�uMy��S��02��2Q�����ޙ�v/
��,u����rv��NT��*AS1����*�̧�����ߊǨ���m/�r�������0�Y�7�^�74�t���R)���d%A����׆�yc_
�W���һ�0ym����y�N�������m���M�G�ܨ��;Ώ4f�)TkgE���,Z��J��ٳ�Ϙ`��e���S�.�7�Qn	A6?|�܃	��g�>-��OJ�G���1�� ��D�E����ژ�׀��\qC2]������ �G�������I�������	>s���P�
��-q���s�+�"�QmXC��]I��g<���8G��Q��*��e�P��q�0M��/pڐK�\�8�= �L�[zp�~dBLj��W9�"�U�O+G���6�� ]���q�� �qa�aYjd)��%��c57|��`C:�'���st��'�iL�w@���vU�"W�v+�'H/�4��|C�Q��i._y�ܥ/)]���K��74#�� ;�RB��������'QːzuɅl�>��:�>b:0��w��{H���3j�0jG���5X�+�j�%'4PWX��|R �U