XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��d��#��wc��p��]�Tz���@DP=�q`k����?��)��E��o��&�U��n���av�4MrLx�y�꠾%y�(��Y�-��b�m�5E 3���#U`�q�He�bɈ�z�'"�#�MbsC���������'i|���S�Ck��Ϋ�8�-j�c�3�h�.c�n����?Z
ܹt�[.P_�Y�j=C~�V7�]0�c�Q.�;�?+��>� NO��z�#S.��~�Hˠ�� �j�B���B��I=�:L��a;ܸ#��~�h�ﾬUK�a��&�������N2x'��O��l��gX͜w=}<_��Ǔ�$�ޢ�F
&,�f)�莉��4����-�
�ɜ̙T,���a
Kd�� 4@G?V(� �,��%����0�J�M�LM*��cf��d� �B5Ʃn�q�AW{N�u���Jc��C���#�I�a��*�6YƟ��=dz#���3�t=��@��ki�:u�Q)\���WV�Zf.��ut���s�{"@���P�
VE�5��;�GP���[�����+S�N�[�	�C�0�zn�m"��ٍ֯|��|E��v���̸rR���.�`
��va��\ a\�d����m~����s�'2��5�i/�.�X?�L��o���G��y��}3P���~m�aSEF���+R��/�β7�F�:&�g�%3�6JL���46���#�`@�M�)��
)&'j����Z�ly�O�J(���Im�"hj<�^����62(�XlxVHYEB    1ea4     920
��T1w�EI>�E��G5I/�?��!6���AĞ~�A�H5P��{���@I`�2�F��@��F$ю�:��]+``{~�	^~���PK��߶��z�)P�[� j	6�%�)d)Os�q���<�Ҏ#�;���\���BL����u!��S�۳�H:��J�uvF����H�^zF�c�GM�:�s�F�\`,���u���j՚�J�4��:����]��A���z�c�ވ0/�c\D��ݟ��G�	(Y?;/� ���tÝ���l͑�7�/9��T+[�{��/�ni1&���I��*_쒐�-%)��G|ȼ�E!�=��@1b��<�.���M|�W��j��fo�o���O�p�eLT��Y��@i�P�Ԅm\�.M��s�cƢ�h�����@*��^�Oޛ!��gO��*�p5���$Y�6[jw��������Vn_���D3�n.S3t��Ī4�i��g��~�f�.+w��d��F^G�7gbl����Y'��Q�1��'+1���̲*�1�u���B�9�P[e�"�+�?c4.)˥�`� �;�N3!�m����
$>�Lȷ~a��}m�J��hC��ޣ�L_b&Y�
@Jjb0�E�D/������7B��.�7�R��?Hnw��YU{:�>w�(v��Jx���3"U�:zK�ݥsتm�w����WD���x�I�G 	_��V4"�b�E�˼2bͅV��D9�B vC��;�`�j��Q*s��iyu�5.�ʞU����ZR�9�"3k�>� �C�!�/����O?n�\u�慺��p �ᙎ��iA��9h,��Vh	`��f�s�C����o�@���+A�/�5-�f	���Zv��d~�'ฝވ5�φ���?-*���{l�W
���s�R�?�`b]��9�T��\�*�*��=]��ٙ,����3��Ң����x���PjS�:*\4�����}�)�
P�p�LG��%��,��pD��,bG���T�����/O�.�i��7:��N�|��^�8�K�c��>��8��͋��'���]��38�_c�qK����G�r⊕ì������1���t縯c�bD*��S,��cunǝ�i�ˡPa����V:�ѩ�!�����z�K��"�O��z:4�2XC|��x��*��錒��n�l�<H��Hx�X �K���y�[�F����a�-~�ܹm���#�48⿽���n�G�{�X�L;�O������N�Z�Q9o����s?�_���61h���w�i���B��=s�yk���������}��P��2!�;,g�m���"ǲB�UV��z��樕՜��5�t2^�/��ۃw:{�v�2l�&��-+��� ����$���7�:NA��x,lJ��5��7(DFO xp
��h�s��誣I��I���+�j՟�z����=`U�}�T�ѵ�-x��f����������
�y�D��qIf���X���d�0��,]k�x+��'��>��[��Gy����ՆKv������P��D#�'��0�x����j+������
���27�?V�B�^;�/y�Z�@�)C�je��q�h4�_ǁ(`<<ī�l�M�l���`��˰{+��=�J���2�W��E� ��=gXs�ͤ;!�@��}Q%$yN�p:BNC����Tr>ֆ�8>5����(V^4��0�%F��x�UW2o�X$t>0q�dR��eU��I�v׿G�'�X'�VE$���m�l(:��@�v�!�U8=�ռ_��x?��OoqZv�^2����yq��#�u���2�������Xs����s��gw�v��i=�.s1
�����:�
��� m�11��WtU�+��� ��K]:�+�D<-��k�GgL�>*�`?d��)c
1GAe� ��l�Z>���rw���ČZ���i��;�0�E*
���U�>��ӄ�q� �V�v�%�7ӻ�yRS��cޜ$w�9���p�A����j"�d�zH�/�uCq{��.:J�Jq��BI�1�Qr������"U����!�����4 ��_�9�hL���	�����e���#��â�>�7f��a��q���Z4,�.Z��Ff��p�3D�}�JE�i7Z��-B����_	���8�?�m��D������v�X!d!���SK�d�ݝ�1͟z3��m��S�U�75@9�o	���;��� %�߻��x����������2HF]Ԝ������a(�i������tj W
�Dv�T?l����%@�iN�=�'���4�qw: