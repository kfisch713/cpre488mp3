XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��'���l��IX��y�@/%�po�w�_��L�-�����F�"9�$��D����ą>��?b��`��Ny�����INdN\�ٗVE�N�ǚ~?��K���d�t���C��E]�L�J.��l�r��-hA��S����xV*/"�Xd�^*u�_Bt�����Q��)�h�Cͳu4��
�h �JmhIhy���[�EtcV��r���x���w���c�%P����߃sN�@.�!yj�i��(�/M��
�i���z�l�B�t��x
�k� �BxP��i��3�!��H��`^-��|qú�N��R3aI���J�l�$H�޵5Z�{e�٭�ᨓ�0���bF0B�l�+ﻔ�S8k���'�'���s��nU���$6�B�>}�
_W��8i���,�Y�[X�z�
"�������	�'�{C�r}if8��#K��!���X� �
}�ޜߓ��v'%�+S:˘!B��v�#?cɃ �?�{i`:EX�!�� hm��������O�ļ�upr�B!�
������G��`0�a�	4��,���cW_ʡZ��2�*�s|�+�R��f���D�c�;DǼH/�O��{���P�UmI�U��8\��V<%n[����)��3�3�2Z�� hQ�t떴Lfn�UGf� `�C��[�^�V@L��A�[�Z�n���ӊ���}�Pl��[��G�c�Z 7<�k�^�'K�!r���W1^��I�K6U�(�������D�C��0��#ŭ.�2:XlxVHYEB    95d3    18d0~�|S'��"�W��|THđ.��5�"5}ͩ�1�<_��2r�믓�G�ꞓ}�8�-�#r���+x��Ӱ��/��2���� �{��+��n�d%�@h�>7!�/H�N/Ga*#������E���\`�Q���؁9�Y�G�ޮ���F�֤1O=���E�	J�	 ��6��U��OM&{�gt��0Xk�߃.|P�U�J����7�O����@L�?*�d���u*؛��D��;�_?#؎l�U�o��Z�gU��V]��|1[��^�7v�.D~�߫'�)u�=��зF�)�">�.詤w$���hm���:ok��ו�7Nr�W�Q=W�&���Ԯ��qZ��t��bm̃�B�.*6�ehU[�m��;�'Q���μ�8���J��pG�?{��'^���ܔ��Џ�(���Ho� wX˷��J�x�Y�}��@�h�@Z5�G[���=�z%)��Ý%���[̽}Ӝf�����cc�O\(s�~�Ҳ�G�C
��h	4χe:%��=��^���p_��)D�¦@ݵ��>Օt@�0g�
+���m�E��H�Aw��,8�f� z��0d�Q\�疔���?D��UQ��"l���/��:{<�Twҹ�2�`�1���s�{�$�|�|?����'H�q�~ �0�8���UM��tv�j�����.;|�e)?U^A{s�����v�%7&��1��_���bX����L���5+�=�MD<�(̼�� c��']���m8#�x��4U�0��/���,��d��$��sD{��{a�uT(����HYn޴�=KwD�^�	��Hc��=`����P+ه��z����2�v [=7��R���X�+�H�DN	i��+iqU��! ����T"v���W:/]�@�m����K�=���]�
+T��fȨ?j"�}��=,1�1WݐV�y�$�r��\�I>Ɗ/�����:��(���z����.��:����Ձљmp��]�j�	�TH�%���jY0��4�z{W�qrϧ���@e,�.�/_ϯP���U���\�kX(��o�ć�%�vȤ#M��G0�z z��LV��=[)���d��3,�~�Z�*��o��V�'�m�G-��d=>>�]�&s�-0/���1����uD,�� lX��� REb�e�X-�'m��ݟ'���Q0)��s�1"�^�x���E��*P�*V-C>o5��-y�YLJ��Q��T�(;&��<�m0�p,�9Ðs�	�a��)��=1��A��`��!���IU23]��P��@j�S��6�mD2��)ܐ�`���:~�(���ZR~�V��k=�ޡ�饯��*�2�r��:�SB�#KYH����m�O������=��Kpd��Z��E����	�|=E��"�QҸ�k��[�c�'0���������e��鸘=x�3G�:�$e�F�������T����3�I)�z����3��rV��!��hC�[��<�h��Ҵ��a�����ԦZCT��L}sLU�D֮���h�ר���W��)�@E{2W���#çB��@�t?e$S/�4љ���4~�t�����o7�Pd��������Jt��d�3nE����54�m8ib�"�B��/��8r����8Y�u�hlh�z-��L�RO
I�a(�h0ٿ����0x]hˊ.4@Yh�C-.����#��.���M�����#��b�jh���M�#���i�B��彛>f᢫����Y��G%���q���U�aX����8a'��O+r~ӵR��+��I�ցӉ^u��)U���_f��/�M4��Dl��dB��0*�����4��kꌍXhBX)�9�{�����J:��\�p����J|�;/�~6+�@Uy��_�HJ����}I@)�����V�u�b��ؗ�9GL��n�38�������5�������f�T����X����.O�֡rY��b�\\.oC:�U!+>{*�j�������܍�-=:���	5��_s�W+��ؠ]r�Ͱ��!˔b���x沞���n.�e$@#�9f7�VY�^t Si~�Cʠ��B�Q��TR�_�����d/���(\w)�p�ѽ��d�9�a�ӗ:�~5Qc�:��S���D�Abn��1�h���%U%������8�tN�� .`��c�Si���x����O(���В�{$���\��4�<ؾb-���!#}>/�瑶�&�z_`m�xT���J�XX��l i��#��_`�Q�`;�iT��� �~�9hP�\y�Q?�2����G֤��-�PV|��ry`cW�ЊH�t�a����Хs[�e��(���ʂ�g�S����$L��4��0A����>�B�R�����>��"�2I��Պ��Rxz���=KFk�����jD:-_��yGEv�����˝�Ro�p�b��5U�c�1p�]���%7�&W�7)����4dW%�X��z� 1�_�݈(C�0�2:���xe{������ۿ�b(�C�P�(��^g o���'�q}u�\���s7K����庋���$�I�E���U4.0$9��V�Yf�d���g.K7K����r;�m�f޺-S���I`S�A ��X�@ζ��>E����$⒍y
����m��R[,�xj��\��x"r��<��!}S�����L{���iQD+���1��)��s4'x\K����Y�� �cHCQl�	9�*iK�g��1��?�Y��zb��L�B
�8�=�˖�U�e>B�j�2�s�*��M�|\4���OZ���=�;Ų�.ħ�������� .��rQׅ{�~�P�m{�а�.3�U�]{�f9RxI1S��|LPq�b����t��Cv��z��cܘT|�����8�����:N;��,�vb��oť��5l ��*J��u���^F��
���vc�HClg�J��gW�E�P7�������W"g��Y�#%�6^߮��$,#T�x_�E�[��_?�I<h��v�T~�+ǉ����(`R(�j@���	E��&F�B5oFb\B�mw(��w�W K���܇�u�� M ٖ��u�����y�tw)�F�=E�`S`��+s.`�0Օ��sXjM�$9��;��b�9�]�� �`���]�`y�����UP1D$dFs3_�hw�u��3���K��k`h�X��]��KO�ڼ�����|!�on,�q��.T�c;�k�{�#t����?��U7����웩*J��_bu����$6��w��`�ڎ!í�n��M:p{�g��<��Y��Jh�R3\ٗ����jI	"o�	\˪�#q9DK����\�,V�Hh��?��v�=Q8�3���T�NM����A�m�Uf�m�L��G�R��W��q�{N|��e�Ġ�ۏ����1�D�Ŕ���I�8��L���!����q��X�Rp�Z�`�����g�Ey����H���?3�]N=s�C6�7��}�AjU x�V���픿Kt�q�`A�u��h9����-#Y���f|A�����럸�9���,3"6�k~��bA�����?x�j\w/�[���Tz�P��_]�p�����5�F����]�CTS|y}�vN`Վ �2oմ��T(�L���� ?�b �FC8ؿ�K�z+e��.U���5���ǃdO�M$=G�u�&��[�G
�Hz�-ms���ZB4q�B4fչ��HJ��Z��Q�Q�ym��:��H'Ӵ�����XD9ųK~f���{�+%Xv�"Н)��CC,{���H�t�8^$�t��`A�f,��a�#sA�Z��ڄ>⮋�e�_�9)���eG�h�E�Rیv&�I�f:S�e�M��ݫ�3N	��Qg�(����LwbCS@���<�?���"?7F��Q���G������-,:%�f��'��q��{�P�X�y��5�"_l�p��;��`�^OZ��?�<�pǔ����ܿ��QU��SC��~�Yx�=���u�n'�ְM|pO�by�:F�������u�c��UA�*X�^_c*A3
	����7����PzŢ���?�<�,��������6�C����k�;�8!q�&&&�(/�8�j0΋} ��tJ����s���1��yElO���j�Җ��/t��4�dJb����H��N
8���E��^�ubU�i��B��=e�����FT�M;�Cd�i�`�I1�b4�'�6!��|b��*��K�?�!eJ쀁af���Z�Y�a��Gc�a	����4�:ÛwK�ҹ��^<�o��K�s�h�)OS��X��oɁig�Kw�@��zdo�8�[����Î��(�u�߮}�u���H��Ҿ� ��k[bLn�Gj��4}-���]�'��L+,v�#���NjL�َ^]���[�SV�xbLZ��s����lWhu��D�����+�b�$LlG���q�k��h��!Kq�d�D��A�/@G��r�bҷCY&.�4�ҁ�>o1���)�������q��AW�t��x����	��7���($O�>��\����t$�FSk+��.�)��	���L{�d�`�{��2��n���8����.�#"�$M��m�T�葷�����]��5�jj<L76�!�F���qk�����g�F�aD�Y�s1{��Z��B�����0(j�LE:����ɵ9��m��-��h�X�>�֋^�ܯ�sY	���>��V-p_N���S�`썺v=;��|{+�x�"y�s�l�q�A��/�� ��%23�`Ϯ5�se�UU�{BrL� Sq������?��r��U��@��c%��3�T�q�]�x�B�v�n�C��\�bom��#R�S������<+�o� �A�!՗o
M�
�&�.k��`d��lG 9(�[0��N�פ@ׅ̇�9�S�]�2{@�ȟ�=)���k�[�1��4K��U3;��
G���pb+��<�5��@��"���l:̅:��������PoU��Y�kB��1�e�O�Z�g�YQ�K�k�Y%�8)�$��#�w.*l�ğ��=��,F�}�/?�
?��F��X�k���"-��ᴃ@���u1WcIK��i,���5���c�	�������#���x�t���f���dS��Q�o��X4�)s��f2���*�be�u� ��{c5�����??�l�a�]�Of*��3k�KIK�+F�=�Ӝ?��o��>z���	�l�L%��\���e`�O��^�N�����������~	u�_�����t�8ݡE�2n�6�<�G$a=�d�Z;�l��T�=,���$���K@Ӿ�v��{̃��g<���MGs����"/  JpIc�g[~.��:}�w��R��6��8�7#�3�P�\g%��I��->���C���۳�|h,lΞRl9"p��l*J߇Ğ�u��X�X�Y�yH�/&�/i�m0	#fE��LpMͰ�K���+���������^��kHe�<C�������W�\����W��bnňf�k!c`��s�J��rC��������%q] ����sVʪ�Ÿ'+n!�J�u̲�G�',���c�Wg&���t���6	v��,�OƟ��^��`�kd�� �����Ӷ���˴F��?�W�=�e4��j�D�|��ٷ&G/yD3�8�1O� ���4�6;�%��0��*�;�fo�EV�)U��z'�s��� �ܬ"*����wQ���*%Ip�7�䰜+�>|}�J��������$N �/ *�Á����}������W	��X�$�7��	PF��O���uլȅQϝ+g`ʥR}�D���0?�0���~��'􏫥(��L���,�Z��
���7˺H��(�	�B�������������)�<֥��Mr-�P�	$�2'd��ayvW(I�
����No�*�̬�2�	dz�c��K)悅��-]��x;�Ъ>����c�����ʛ�k9��4�-��Ulx��-9,T��r&���|�-�|]�eP6����f��9o���G�g�=���	���O����(�֏�Թ�P
�Ls4s�u���V=0"�0C��53����m	�ls�ʒ�8B����1��mI�in�!S����3rwED�����a�ݠ��{^�.O�8�z?��YO뛛��Aȟ-��'�7R�ʼ���%J�N�̉�Xr % �߼�Gp��