XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����i �uV�n9�Yﯴ�W�]JY�t`��3[��c���1���!&�'��[�����f�䟧)�X��Ñ=�/ �4IY�)�trS��Y��r��<�I��]��
|��p|��ؼz�3�T�TS7o���2��w�4�˭�,�^���Rv8�/ז��4���&�c�YT&iu\b%�3e�R�� !`�]g�z��Α��\�V��s�|"�N�*��Q��I�^����^�Q{w3���Z��}nU!0���Ve	���oW�n4n��,F~�s)�L���;`�6��-��.e`8��� Y�g���.+vl��U��_��4�\p���u�#�v��5�L[8
�ݐ��Ψ��{�+�hkE��޻���ڀ���`]��S�$����V{� -_>���;�A�v�m��l:@��og� �s2�$�����F�/�-,ҵ�d��Ya��	�"6��?٥�˯��@f�<c�t^f�!Y�C�	��Y�B0��'
���(�4糖�o=�&h�&�/w�ݔ��Q��2��MO��~�TSߒ�j4�77[�w��C���V�c�a��r���^�Ryw6/d�/�~*�"�`��X�=�}�ԐE�21($'V[X�b��N�wm3\w�j�ߑߒ��]�{v����؎|7�8����h���7�qC�.SR���Zx�������m��h��x-,�>UVW��u��ݚ?=�H���Ef'����f�iǻ����-��o-��S7�хQW�ShM#������̉&��QXlxVHYEB    5d54    14e0nvh��`Id��d���As=��k}CX�F��Z�;�\c��ь���`4�ᕄ�ޜ�`���ER�I��!z�򣫳����]]w8�`�@��i>�L�?=Z��F@T��P�d������^�<��o���%&�/h?d"�<�y���2FF�>°g��S�iú�jG���$�1��\�ӣ-]������S�eY"��x�*����Ȭ徍����>nT�b���ކRox�k�B�'�/�qu�T1�i��:zJ"�a����5&aƺaPA/0>��j����3R��Q�������~��A_����A��z�b-y����`_&M���R�-O� xE7V�@ȍ�i��l��B�;,f�g>x��
h0�Y6fy`���&85?��A�</oy�������W�����#*B�I�6JŹ���� 
�9�� ���]sQ�1�ځo� �H
��ڂ�6O'�"��C`�f�(N �3mc_�a�t�*�ph���(�S$/���B�K�=yE�"iI�a���S�|���,��;j���*y� �$��7F�Ebu���<$m�������v	�t�{���^#�N��ȩ��jg��A������6)�����#��a��Svz�dN�)��7;1��/z��F+����\U w��y������0&N
�)�6��Eg��)f�k���ƞ�eH��Y�o&��G��$������_  �"��f��|t��T��K�7���B������7��N�S���X(1��^_��#{צe�F���^�t�T�G�kI3��w
 @�/�!�c�C������M�w�[�X��N!�.�q�5v$11�5+�@��#}S>���;KO��l<6E�p���c0�����f�����g���6����p{W�0��A��(���T5u�F�፝H$�~fװ��'�ˣ�D3���{O�U�x$�8��r_�B�A�Z_��Vb�H�6�gȧ9�lon��yJ��
�#ミ��U����v�D�|!5�@h�\��~��G#�%�i���,e��s� ^�it�(>����h�P�;޸��,�����h��N�,���z���pk�
��0D����hYط���B�b�>�C��&E\�`�T=���������J
e��`N�"t��\��ʀ���H.?�*+��g�. #0��i���ep�R<�fh�����w�d���u!��?{�͢gg��u�k�*L|�X���R�4ڽ|�:���<p�CSǌ8%5�7�1�5�g�/6�3��'0�i����U�Z��Ty+3��)h���T��{2`�R���1�����+�d��3��l�
W%
/m�0�P�Q��6��8��f$�� �u���V%�ĸ��`�Դ{F�(�q�z� ��`�ud%�]��cyc�U��e�5/�J�t�ߡ>� ��豴�u��v�+�q]������?��T�v��'�4:0�[������-g����VcV#�K��0�������p�6&��
ƴP0#Ǆ�Y�G�n���0�\��$�5L�U11�"��!�o�q�d�j�zJi�K8��^>� �+�H�c�
�,�S`~�oc�s%�`�.��mǓz�$O��kj���Do�O){�0l�@O�q���R̳�,��8c��~+�|-Y/C#���_�������n_.�}����.��;��Yrq���U�Y�X�ˆ�D-S�ɈT�w:6�<��m��2$�ޚD��\�wH9I���5��8��.�^Σ<)�E�D�6`�f��]1��{+D�m(Nq/�Z	�6R���j���D���)nY�Qz\����@#%�!�����s҅m�_Q��9uΛ��'hS|�0 �,�^/U�>�Pq��+�~1��z5�8��Xfk���.]�_x*	�Sl�Y�U�ߡZ��֖���ʹ�)BtR�y�:u��nܾ\����)P���8Q���gv{Z���%э��>�?���c���oi(BL�Lt�_G�
�S�[u�ے��ݶ&���PrcQ��I;�0�C�4��r��{�u����˱�e4����urƢ��:��?��u���yD�q��'@h-���"ܞ��;��������^S+9L�_�ޙ+��8�`G�7A�Ր�����	y�]Ĥˋ2y�OD���\��L�q��y��И���=�-��(��H�K��s��"l����+�}r�Ŕ�-�8�q,.�Ӵ�3��_	�y����ks�cʽ��������n��ON���m�����/Qp���4�e�� Ռl�GΛhC�c���hb�4ۭ���$<���5�!#e
O"�w~�A�p���Ed��:o��G�$�'n�0�]&�ea���s�ZY�z���m�E!bKy�&gtx�ԉ����u2̛ЌH���C��#<�����l�\�I,�{y�c���&i�5��ny�Kw�F�X'~�� �"�B/F����`�^ג�
�j��Xz;	�����&޲˱�cv�`�'���uS����G��C�x)j\�M1��iy|�,t�]k|� �9Uȇ���r[M���S�2�|�"{�<<6�U��ё��
��8ŝLe�Z���ɱ��nG�?*��/ܚ}��o�#x���_JԗrPZq�ɞ�i��I�A-�d�EK��O|T�������E��\����3<	*��E�w�C�xQY����H��3ՙA�[[��|�(%�+1��>��x�h�� @�+*.�m,gV�ķʏz�>ǭ�t�0�<Cz>T���ib��?�R���l�A�/�ށn�Ue���Z�-�Ҫ�����L���0�0`{4��yb��0�@o Պ4�|[o�J돪�L�egC8��r͹xB�jQ&��(!tP���V&��!/�GZ��Qf�i�[{~������ܐV�Xg��c��w{ 82�1HӨ����QI�I��5g�f�g��W��S�4s�V�&Ӕ��((f"NL�9\O�+R帯��[�8���y��A�L/G�);6�v�4���I�y3]R$���7� ��ͪg႟зԍ���z*wE\JJ��y��â��Ď*MQ��R�񪃤�z����!���l�;� �t��Fb�1��h+��@�"�`&$!�l˲�xO3A�>)�1�c�!Z��8�����t�&~N=)�Bq�vfh�i����t�f"4yg4
�ac+a�,<��S](g��& �"�se�KF���2���|����GmB�LBA�$�+�-&�Ht�.�"%h������ ����֝r�>�I�k[՚É��0|lN���F�D��gMh�`03�߯EuT�9�W�t�LSp�#���o=�u�a�$R���o�O��]���� ��^�Mu��w):��H�����"�V���&�[���+]�(F���(	�g�q�jCw�ч�]؜ڪ��W��<֟�K���S}EK�Q��^�r2��F�C �6�&9���P���G���Zo�q>=��L�G\�4�G��Q��I���E���*�j r��I9���R��.�T�1Ţ+� X��2%�1�a݆�vX�����Ǡ�Ɯ��e�L���x4Bԃ���>I���+y
	 n�k�I	Kߡti��ZY!���Ձ����Z��� �
̟��q/8ϻ|C�CQ�P�~�qv��ۗ0\�~9�17;�Q4g��v©��^[�ڵ$CI�d��e�,|ܬ���D�3��2I��D�"��)Ț.@l�{�+	�m[j�~��D�@��UΌ����'�46�[��JC�c�Q���7���l��@z��V���� ߤ��С�k��?�9�~C�Ze�m
�����RG�[T�J{��d�s�e��IDF���U>��ȱ�)���7?��/<�B�����Ű͆���x��9#ʊփ��GqC2e��X>��,ݥ;mS�CAڻCT��&\HA����Q��Z�d�;ٯV��W<�@�mE�=�0� )L�@:��l�?Kӫ�|O8c��u
�z��E@�LZ�Q�Ut�T�_똵�z��\Le]�t,�av�0�k�6 ���T�[�w{'(zt~g�'Θvq!eu�k��آ�����}���5Ջ�f�&Y�hO��s���b��Ї�A,�&�Ý] }��yY���e;��S����"D쿥l�㒂�H��>�̌�C�<ۍ���[^��>�Z���Y���a�%bm�3h�����[ۊ�>�w9١�G����-Q5$�_�g�� X�8冚1�:nz����;zB;7�J��_T }�F�����l�AV;�3�"�4�4B+S��sxб|�]��5p�+z�DZ�X6_�Ǜe7po�{�ډ����r����<�o�q �xU�s�,N�߁�	�X%#�I�l�c����'�#!���8��RĬ���� uU%���(�(�u[3���_�4'M��T&�Zj�D:��&�6C@=|��1���\�2�l~v�ye�G��V�E�r�:��r�K�V79���#�����7;�YѬ,�dn�E�3��29���p ��$��|_�����VDx�d�h�ORҦ����.Of3�Jۥm�q*�J�΂N;���N&�O!�yJHr�s���f	�~��~��Ҙj�Ptn�(��.�	.���C�����r�V뫩�g����=�� ��%�$�*{�zE�v���R _�5,�"�\��G��#��Ir!��b��3�U��l� c�9Ȃ��Ij f�G����J&u����V$��)���2W���G6*r|t!0�|��K��7E�������o^��V��� s������s�sQ-H���ͥ[��%ALgv@�`����,i�6���s5����#�><���T�2NQH:����:���]�B���˝)[�Z���8���c��+��OZ�h�tp.[���q0�C-y�����P��|�2U������9�S�w��;`�BnR���Y'H���K~F���+���?r�O�HrX�=\���u�{���+}q13�x�is�2��|�x5��X���[���U�݇��H����\-���6q6I�R'g�@2<��1a]�īp��ү��<ܴ�Ђ暯�]!��NØLd��_�tE��5'��f!W�%GiA��bպ�7P��릲X�j�<ɂ�/�r�����\���6w��j���7�zk_�r��ԟY��|�����]p�V&����]�2���r�:�L\�D�/�3l��P�g�ǎ��'pk�r��ߢ�5������&��T�Y�zW6<
5	��>�T�Z*y]�L�"��C#��W�Cz88��