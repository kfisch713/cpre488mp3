XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��?+�&�]�va�WB&'g��a��_v����Zi�O�Y�y"0A�Fɋ׃7CI�i���K�EW���VwGa�� ����B���4��HXMR�[s�vU	ҷ�4)E4Ɍ`�<�74հ��{}X��m�)!Nu�v]�}��Ke!�z��������#�:ǌ$f� ^8T5�B��^���S����7��2��ȁ�]{���_?K�|�+�� Sp��$��B�uyo��r�è|r�N�q��ߘ��v�	PN~s|� �-����-��/I��5Ir��x��*bP�j���|E=�ێ�m�ɜ��Ѓ �PG��ą��R��Nt�Е�Ե��M.��"�^��!7���|�P�s���r�]X'�.���,�)uZst�)i8Ǯ���t����lPT�>Kd���ķڍ�	kt6��\���`7fu}���:�ѐ���m������D/���Й�Dpb]�G\+��� ����0���!I� ���u�+�_�u�2����o7��vù�X���{�F����bg$�)Z��Nnw�*|i;�����GG�li�ҏ��i�y�',�b+[Y��P������T ���; Ư�5�c�h"���<R�z���M�}�</p�֦J̈́GN�\&ɨ��f��}�GID,xE[M�/(!n�n;��|�WՁ�r��\��5��_I{�d�v_s�#ޏk�Ħ`�B��~(͔_͠�*���J<sp�P��n����?
�8[�������V�>��XlxVHYEB    82c3    1970�9��B"����BO��p�*���=�P�!�S�l�yՖ!��m��A��2�T�E�@^���R��M�q�at�6�i�ē9�[�(-c�qvgÈ26�E�|*ǹ*eB5J��k�����':ѳ=5�k�j���$F��. ?U�#[u��U; ���$-����U��h��r�֔L�ѠMRJ[�Sr�_�_�]ܳ�̗�f�G����$��6[�fb���U(����ܞ��N�n�C�S����l���d���� Qݛ?F��#7{h�m��Er{u�V触��{ܠ*��]�X�oE�C Q�57\��)�@q�p�2�IjqяX`��K(�DЄYy��6���,�V�'�uUYGT��#�A�rT��MZi]��;��O C�I@D�Z�l]1�A/��{b�ش@�u`�ԫ!�b##`�:�5�HZ-��͎LA4Qf��ˀ!�b=-�����z��1<m�k�� )v��9���\�dL������{9~�q�FK�ͷ�� n��i$�z�.��\h�G�?'�y��6b�Yl�{�!���Ri��~u���)��WQ�O&��yj(\ʛ6����̈́�@K�Q�3눽����"�b��.�i�>���i�Co��xj�&7���v��̐�z{U*О���5��O�-?�hӛ!���:��ZcŃx�
�o$��åi)T�lK�B�1<��T�L5���2dT�H0�}�^�ľX_��[QFɛ�7�J�}��	�7�ar�fb�*hB�{�������O�}Fh����;���9�-�#h�2m�.�;�����\�}�����"�}eo$h�9�U۱�5�+����v�i�����-�	�-�(�ރwW���3�
��/}5�{��KZ(c���:��f����L���j�KP&l�W�`�l�$���>yp�V���Cry���?YΙZһ%������:��TGfc�sB`M��>W���Ҩ�g���B~����M���c�n�g�W%�1�ȱ�j�"��v�v&�R	"�I�z�C�ԇ773�Y���i�WW��w�@���I���9R��t°l�����@��dH�R�C��h��?.�Sd�YI	����^�NS2��.8��I��� �P�?/SC�2��
�<������Z�q#�����4&�~]|S�a1�`��)���zUb�"�:�/#t�*�AM�>������0;v��X��3ϧz�`���ƽ���8K7+W^�
w���a�./�co�j�z�浄I�?O���}**��BW+��R�U��p�Xwڒ<�d�<�+�%�Zl�0�-��B���TŵH�H
��rN��*���x�K�@ܕ�BK�n�!�K��>r�6 E���!]"h�������6�'���{ɻho��hҨ^�;�%�`�M&��4�y[I�|�^������n]��vU���#��ZGQVp������� �<* �;�%���ԊQ�Txm엙=-�x`�����A�����σ�f~����2|RۀK\��l>����u���qX5��£����R�K��ꐬ@+��v�<cB��`�'��e1�W4RH�ʞk]�w$:����!�|,@�.1L��lO}�M䇮I���vn���uq�N��9����S�S&�k�Z���ٮ�#VmO�lq@�4	�o�O����hj�;�� �̛R_�`T<n]��(�rF҃(;9�:3+@g>���Y}�Y��l�v�>G�P�ɨ�c�i��~��x������4�����K$Ӆ�CթQqG`� ��NtT��\ �vZG'+�bBq}��&�-�|@�N��V��{#��+�M��p�������^�E:��p�4xY�e�wrt�j>�m�����g{����I?��hz?�.�y�t��I2�xX�����G�]cr����ՍR�w"�2�E�1���mZ�>�IWܡ]u��y���7{��f߂��GH5+~��U��оԭq����=ί��Iw%��J_h�!3�>cá�ӨS�����Ԝ.����C�C��W�܀�$m?�-��vM��:Q�ׇb|*H�NNzKI�ZR	�aȞr���Z)%f(\L�� ��I"f�vv>E�O��w��y�G��u��r��n�~=P������%%���b�n��{)����N�?z��>�o�_�O�+�M�ߴ����5E4����gx�W?C�@3��N��Q�1~�R�����ޜ�X��!Sn�Q'\��n.��b.���b�MN{��).ƶx [�QM�Q�{�C+��]�W�`��Í��M�]�� �e��/�Jp��7�y(������Fj���BM�7?+��6Bs��7�8
b�e�3�<y�~VD7�g�muO�K$�n}2h �� x)>�Z*��R,�D���'I��Le�bA��vn��R�?�ig��OZ�\�H�J� �#��!��,�/������6Iv�V�[���	���X�m��#Ƒ��g�������6FR����{X�FE��ا��U�ޡ��g�K�f��y̾�_t���o�8�J��y�yK��w;p$���uYLv�Ep��Xo��H�|	��za�+/��b�6�\RyD��aB����(����l�|[1�7*{��J�X�+�����޷��yT��	�C.C�l�xƕ�M�t~Yn�r�8b7	X�_وmBC�����c?�L335�l]�U`�����R&�S.f:�1�v� 
�q=f�&mo��Q��~4:\&�6;�Z�#�?�] ������iv'k��4)�YY�$w�M!WR��o�UE����p�����.Uj�6f�����f��zzaδ`\���QU�-�h)��xՈl2�;�ĴN�k���:S=]y���k��Q��U'���~h��3ۘ~���,� ��R5H�?�eg�\�ht��BoW���h	�;��p-I�rǧ���TT�KV�='/It�68�G�m��\�~�\��q0��c���鼐Ծ�	g���Wff�z�J�f�{�9#}��$[40}eE��iJ��:xN�g��� ������Yhz�Q�ȴ��-�Q��XY�D~�b
�:r[�m<�육0��Ʒ���3A}�~�#�`f�F�P����uGQ����}śY�I_}�_(�X�4�U�}�^v�[�X���b��8��0����o'�rZy��3�Yǃ��ڣ���`DvZ⦒;�%J����*�R�j��/��b蹅��T�ч~Δ�� ?ȺwҮ��圝�@1�=u �Rh;u�%��K�%7�n�~�j�N��qm��lD3��-m��E/'�>ʶ��ʩU����5<zY����q����$�;���h�]��JF;�R�7�:ݬ����fM�2�F:�_���ld&H�Ј�������w/��ZJP`>�ya��V����W�?-O��	���c�D76����,��z���D4���i[:kSK^I#|XP�h�5���L�IR��24�Ap�N��w�2|g���.�6�?��!g����:�I�����=�Z��L�+���#��T�7NZ��7u�|'���`͑VE�ZE�U��q�Uo�ĳ_86�t��#���LBM�hT��"�a,#-\���8��Y\��>���r= �ƙ`���ǵ�<zV�����KPK\�G��97�IЄz�}�����?��{�.(���h��:0�: ܁�j8>Wi_��];����$0kf��J$�\F�Ͻ�-���6(
��#�:�<�s�c� R�v�)�hvR�/��5�,'��B�+�h�w�7���� h:��3rj�hH=m�\GK�E���8'U�څ���a aڕ�������#?�fq2-kߵ��D�NB�G�:aC���2`�Z$�\O���/bOK�n�~�Xz��f05:M�v�'TGL����`L��?�FX���n��H��^�7��F|��L6]��c����]�d�Ż�`AQe�׸�]?�i�ry�R&�t:�B�"�~Ez���ķQog�&��%^��l������4���ڿuٿ؀8�]��`�ʬ$��$�#�^Zi^^�8d��AU�+ќ�o�T�	��5�B��G
j?daj��U-zY�c\������Z>L8*��Fn���W���E,�|��!;6�Rd�����8�$S��\��z��Q��W�8�^<��O�N��`�g�-�O^�P7�㫽��	���b��"�bG	���i��ޓ���ڑG�-�X��4YN����­X���H�I�����g����ķҧ�_��=�R "�W���/Y���r�����յV�V���{�r�k1��M �!sW�օ��p�O��n�>���|��k#.�$m��[0n�)���s��c�V�i���<�������A���<��0���bi�8G��}�⾒]�$�|9R�6���� $��(gf�iJ��}�,q#W��F�e�؊���qFAM�4fPO�7#8�9@(_P?O�Lr=ƧrJNtj��8��{�ppA�Cv$���B�3hQvPJ���U�n&��I�xAK�8���	?��q���皺X�.��/�4���cj�Ӌ$^`�,M��w�=�%�n�����1j�����4�K���[�Nתy*	�����˩���:m8�\�$A�ixA^��?0}��R`W��im��Js�C�y�驏���ڶ�k��\��D� m[�V{>�R��\�h�ХA���T��JN�ʪ����b����C�̨c�[(Q�mi��ѾR==�-6/u���)s��:�9{��R���Ւ��SMI�@�LJʲ��\@"���l�c����O�����<��)͒�������PF���7eN%�s���sb�Є��@�;���J�N�>J>?����q3���q�D�A礼�=?��\)���hjRhЃ�SA��o�G9!~�~-�VFiƜ�u�5�⬲$��_�&�㶣�W Ii�OU\e����E?5ov�$ˠ;!;��2�8=6����^��Y��o]H~ن�Z��q!ؚ��7o��T��A�����h���m��e�ܟ*�q%�4��	�p�|�V(Q��u�-}L���*Y����n�P�	�������W�����o?�K`�`��2U��:�$���t6Ƿr�#��r?`�RIؼ��CA�Ah'm�j������or�m�ڞ�Cc����"�.V|���tݽ��,ٝ
���5�n��I�0K�r���JU��A"U-|� �5H��{7���W�:�55�6�1V��kۏ���W@��H��j:wa���ƈJd�3�on�:ߍX	h��`�Fs<�"eW���b�_��v��V��v�Ia8��f��͎��aN�E�a@%
��:�(��-c/�������O�D�U0++�+wc�k�\UB���)��Xż�iQ��&�|v����@����Y�@�����c�#��L���Y�=E>k6�]j$�9q\(��4�X*�i~��=G�R�3鶜��Htg���u���ĥ�~���[��l_0��km����"�v������� ����S��_�>�8~5���LP��|��QG�-����R�r�,�IwEh�ǥZ	�d�������'��z�n�m�Ki��w�����&w*{��#�9B����b��O���������vK���7��M�B��|k��p�飸����z.{�B�~VK2d��FY<�dl��A;��������Bs��Wb}�V3��Д� .���ޯ�Gg�(˓2�ҙ�Qo�i����î�ȱ��좡N�\�Avg�1A��K��zP��=��{w��f��h;�Pt�2vMH=t�`IZMX{ �ǐV�7Z��y3�9v�hvw�=��H��B���`�!�8����U	ʄH~�u���gbnyW�c���漖���ag��:s�Vm�������H?���;)����cZ�~|�Vmb��iM�mr3��:��a'����:r�p1J@#�&���p����� (��\9�'��C�*"���.`��Q���Rt�}Hk����qA�cY2�+~�3��b֏1��kjUo g;�l��?��QU�a�F�Ԩ��V:��JCy�|��؊A��
e���զ��"��.�f����,�P�ӹ_/�q���N�u)�.�<nƲ�����^��W��ןϮ�VA
��~v0�������A<��;�cp�P0���v��D�I3�{ 1��휢p�D*�Ek?����U��e�-��A�>	|��w"qΛy~]F��w��s�G�ya����3@�8�wv�|�|�]���M��b�ئ��=�\=Hm����εKL��U�z'�a�t2�?�V0�
��K0�F ���;���_1��Y�X5N�ZN�YD�~�B�z]�>��# ���>�@�*