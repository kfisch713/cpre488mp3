XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��'��f�+g8���깍����z�T̉�&SS�7c6�s`$�Y��U����P����a+.\�����~���LG�������L��ȝ�	���3�W����ť�'�G-D��������N╇9.���NI���	|��\7;�A�X�*���QIoF�U�&�Ǥ^u��-1ߍ�L�f�q�	���y���9ڷa��Q;UK��N^!�APaű֌j�\L�!��!{��n�f�0d��jt�4_��{+G�����[<*��$<a�Q�="����my�K̎+�D����,�&Y���O%��\�>�B��ʿ\c�m�����r@z;ljC������3��@w��ښ�����MZp�6o����{���̢ޛ��ڔ�W9������jBmP��o�hu�lP��>~�?�!�� �_q�����++KI!L�O�g��3|hE���$��4�q�STg��߷o&����,� �d�k��}�X\ *݂�[��q�a,�/F�_�'iU?��nE��<��<N����x!s��B�~�Ł��m�H[lK�g��1U��O�L���ٜ�u��w2R� �����+ѭ �Fl�M�9��G
U^^�;��G8���t���X�0�jlSo�9y��1}��"\e �pR��6��h�]]��ҧR6�xK�Z�J������8�Ϻp1�������8@�j��{�R�6�}���Ύ&U��G[J�.J4�6�V�P���c�F�6��W�
�9�8��a� }!��G>0�z�;XlxVHYEB    3c24     fe0�>.`T��!�վ2��,M�pg��i�ܢ�#2Y����r.h����qyX��������nV�P\->(���Js?@�m�:����;�9��4rd�_�V�kO�"=�I$��h��\�
|�Pk ��!�E]Ճ���<b OZ!��(��V�+��)�����'m��p�l'���J�ȈoL�b�I��%4���G��$i��%`2^!��ĕ�.������ڻ���DI�����CD9�%�����.j4Iǌ!���G�-�n�3�?��}�x�N�y�	��<�y��w�ߊ�` (����Zz��q`�ٽT�3���7��'����mb\��m��hܯ ^N�p��2�F�zt��Ц�u���e�	��4w�"繋��̷� �,Oe+�[�ܜ�+��X�����+Y���t�&G�,�_˦~APʴF5�I�[K����2plc^�`�%t/0�������I�A!p!�3�gm���D��� �ұ��fF"ER��M�z%�����sy�O��l��O-��5h��Z�x�T]XIY��lw�) r@};��C�8��WA!r�(��7������o8��r���6'D�㵞gf�紣�;O�Y�,���n�#NF��a�Sv��9x�"���{�i	b��B��}4&���%�6�sb����>�d��=�^5[ș���)�gl��B�\$z�/Q���Cc:=t#ɮp$h�b�e�̓oIch)A�	�  �|E��?q]��K��D�b[2�m8Y[�[�B�F|��z�,o3���l��3.���b�@%���,(.b��ް?��$B������mհ��h��$�1:	���h����{KY3{<��|O�8)��J���B���Fz�:�� G����o�n��$��!�2�j��ۼǖ����U��A��*=gl��"��_�?	�|��}ې�j9�Z� �/2���r�%�O-��Z�gX������Q5��c���VA�:��K$���s���?�-1���+�E�@�>[1"�p��+PS/���J�{��h��,�N�4��9��`����ϝr�,rL9�:n����$��8�6�сyf�l;r���u�$|o4
x�l3:B�@(�/BF�o�L��0<�)$�#k)P�2d,��=3�ucdc�Orwy�
����IJg
�4�	T�{�rD�M���O$m��k�8��<&F88��Q˞���Q��Mg��p0^��?�u~6�̍���ˋ:·���BJ�q�	ܺ�9�CEt�7���m�`�����,�*ׇNs�����A��K���Rm��I�Ą���!&��6�K2-|���P���44ɢ[j�oU7#O"�܎��N�#t��z�Gx��a�e��>�v��9ƨ���w�#p5��üg�T�2����;���?�lz�"��!l�+�:�W�3���WMo�7�f$�#.��H]oܱx,0�L42,�Ә�u�[����	ip��j���c*j�C|޸	v+PH ~N*��q��j H�so�$>f�aM,A��i���s1� ^qG^�
������q���VS</t��4WǑ���\Ɗ�XI���@���S�NK_��>������_��t�ȣ�H81��QѲr��R���`���?�B2���(F����*/e�+��C&�x�VmĔ�y�-��B��qg�VUDz�LO��0����Qӯ��ux*tz��X���f��Sp����Cr���6�K�d�[yt���AXj��E������kvB\V�[�VBVJ�9Y�C�ϻ�\q^&�j��|��i5��a�-�>��c�e�`��XK��'hŢ����;m�X^�~Nk>�v��������ML�u�>Rp������f�u�fD��{l�X��x�	ܨS�P	��ʻ�ӿhrUgz����:7�0K���»~�f<7���� H���m>�N�
��T�����כ�8�v(�~�NG�B�I2�(�S�G��������'��f�ٝ�A���Y��ux[�+���L�1�����n���g�}NjE�vy��WG��w�UU����)? ; b���ňĢ�@�E���ot�yF{���5@�I~���t�B�@J(B�a�ld���/T�ek��\�Q�';`o�]���]��=�A�腛�؏��b�7V����$��H�(�S�Ȭ%p!�i�q�8Y5��x����:�C���+[�1˵�W^�K��E�U�5��!��4q�F���F=���}栜� �$ʲM8ҹ��$�Y���P��A��OM>�Nk2�#yS+�)�>o��DB ��*�k���� ����6Pșa����Jo��
��ET���U�#�4��]h�ij��Q���g�%��\f��Z�&�,���aʱ��ϖ�:�1VV��c,{�8�����,�V�������=�Q�c���'�&�yK�Z@���v�����7A������(O�� l�V[��.�ct�i�a�4���:;T��1�y��~�0�\�q��k�#�Pia� 5-�zg���=�2I?���σ�����5���2�T��}��G��6`�JnỤ}�4�`�W�)�G������O�t�����=H���xny�]Y������*���`M���a/ScĩC]�$�~SF,�n�|g�׾���8V~��b:��ts9�K(������n`�hD��}��/���e�)��#�O]����Q:BD��l?�"�
ڸ1�U�:J�OJ��/'��9�S��V�g�x˕��mrx��O��
��U��0�����_���O��YfNGp��7��ɻ�L������޴9E�t�.4ٟ,K������4�0�VϺ~Z�C� ��;w��E,���bP������s� *L��8�00�O��H��Ё �)�FЉ�6M���|�'�NN2����{1㭄��fԄ,J���T�=��w_������{/5i�Xr�x����B�\�V��Z�e���*/�B��?�T$�T�W�.!X�-7]��$�a*eYo��7���b���:�������H} )�!ib�>����e��q��T�zĪ�qs�	W�;��
��]#�6�K,f��/�_d��']�6��dcrε�*���4(V�`�,�^�wᇘ�Qk�DĠ��0k. �6����M�o�����dƹ]�q��! jAF �S�����lk"ZD�=E����.6�,ad3�r�X�� ,�+���q���S�."a��qfT�
uA���L�����"�BE|Ы�=ڴY�bROa��a� 3�8m(������"&8oI� =Ѿ߶-�m�l��[���vHB�~�0�um���2qnEZ�d,Ak7�}R�-�/)<D�ͬ�l�L�uŌ!�MA�S1	&����P*�(��2�ȱˋw�T�[��>X���.]�֤�r���OOA�;zS�0�]^�����P�L�zy�-�Cnb�G���1�!�sv�ە�I���@F3�#�Z�{����ՙ�G,P��M1�T?����X���LC����M}�Ƣ�����5C�Cj���`�Fa�H�6!64�a��� ��a���PŨ��K�-AЬ��fl�X�dI9B��fL��o�f�Wy@����نuE�uC"Z��/�`?~��]��"8O&9L�#qB�>->�|��pH��dkY�_�ƫc���w�[D�ZJ�5w 5�+�m���wQ�{���+�d���GN<3�	h����L��ప!�~#���>u@�
,�!ë�;�s؁���fZ�_��u��>���K�H����j��&t��� aVM1d���e޺ o����� �.�֬85d/%V
M�����m�4��/Qq����o�Ӓ���m��A�腏�
]~>`"Rԙ��`\n 	����u��DP��db"��x��XW��_tz?ܘ��(f�xU��qzoG:%9+�vi�4Rڄ~,��
�噱V�n
W�&Q�O�\@oId��j��g�� y�Gc�����