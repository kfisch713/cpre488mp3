XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���ʞ^���2ܭ�|������K!y����@�W�W\���g"�G$���Ї�n�rT6h�!�G���(���������U�~��iO��Qd��9�՝��S�6�s@p�!ꖾ�֠�\<�l51��v����cH�Q�|��xp���^�1�.|j���J_ ��9ۖj2�A�DN�lt��xY��+�61j������x�14RG:4�׮���T����0�HJJ	����;IUŢ$�?�L2�=�^��Id#��J�H*%a	��ߎA�ͭU�ߋE�2LP@w=�4"z�R�e$�����Ϫ>�K"�
���P"������wԣkj�c||�z�u�W�C�$��gkÆ�A�#�5�Q�Nbf����.{h�	�	
Y*���Ο�k6�$�%ꝧ_VZj��9U��ԯV��`�6��q���J"�>��O�A�[TκwGKqe�e�r���G�����~V/�Ҧ�6s ���?���ܭ �] )�6��S�<Bp��P��I
��Y�#CN���Ȑz��E��c� ���}�e���[|�[�9?#sa��/�K�G�7�Fx�ú�Kt���06Ƞ��}QWcP��
\�������l5�UU+|ޖ4�2*w�b����0,DC!4���c=p�D+t�� ũ�i�J�6(�����B���_r�e3��?ʋ}uB~z�F�|U1��!��+�@��	�/f���%����ii:��"����L�#���P�NXlxVHYEB    4b2a    12e0����[�!�I�w!�N7��Ro<H��ӓ9h�dO��a��8�w���\�P��iԘΟ4���J�ŤȬD��.+��9wl�j �X��E��`�3��hxG�8���)AtJ�6�Uϖ�h���Q#[���;��t->#�1-���q>�L�I�'�v {6M{ͩV*�]�֑dp�A��%-�!Hi@��6~�6~*⏎�c�5-_B�%��=$�h�����ӞUV��qf��(%������K�N��d+�ʎVh�Ð�i륉W�x��|^�ʰDy�5���U+a�L�����^ۨ� �P��^��a~��f=	p�{������l��:��:zHR��.��8����q]���=�'��_�/6�����K\)oR$-�qinɏ���V�~T�s{�^�eDVK#ӭV�rf���8�=pZ(\�ʀ�zُ-�b`���HM'cnsP���|��p�fCI�'�6�j&6���C�Ƒ4N$}Um]GU��%���<h���ņfo�&#����s��������\^+A�?��j�˭�{h��2n�@�U��{5�b"
��R��ɥŰ�=�(C��<��2�~�'Su�����v���ǳͩT�Ɲ ��d���O�0b��5ǙVG�����ʧA�8pg!L�����B���o�뺥Z��u�.�mO/��_�O�㜓�) M+�,8�w�|�k��EM7��o�70��d�b�ǚ�����[k����n�������ye�ܢ����9���nL���mg#3Eʵ�Lh�lz���X�֔a��*ZN�
��*b.�A�ִ�;g��.�Aʝ+�M�KeF!��@�&Cy��Z��n�l�4e◨�p��T:���hS9�^kQv^5��xB�4xC�
�g#����Ď�d�$p=��\!e�?���#m��*Dg#��Hfa�V��vQd��J����d��f���ìDݡ]����<��Dβ'��@F�|mS��*_��-��E��2��ԇ��'�t�>F"X������'Ŀ�7\���Ƣ�9]1=�WәE�Z2d��c�-b��P��E��ЫŁ���r
-u5�$n2�r�}��1�𷭹|0�I�;��빃�?�.G�O�-��.5"n�MH���-Y{�+�(k�Ό��n��R2
noǝ����~�;g^�S��ēs���&̀d��C��J�V|��%���.ܜ��}۔s&(�c��2!�8���z�Gy�w�E_�/��0&�m���vV�6�H��AWr��k���$3U@�ǖ�YLnc�ѵ�N��R^Q����i�@P�V1=���"lC��8�Oq��e�#�������"��>���#C��wQ��l[��FU��"p.Ɏ�>�jpg���N&׮�Ĺ��1!Cu��k��Dfm�ߏ������,9d���br������^��0-aE]P77<N�c�	����3f�s���s?ߠsZ:5��l�r���ԞA��i�]�m�����"/��ݻ,i��	kDd���`��η8l^jx�jT�{ �`czS�G�Z"'eBO&��:�l�I�<�7�'�p񩐍$&�-[���i�YM�n�B��ͻ����A=��k�;8i��-$	�7lS�N0'���syT�n�-��H-�8��N���	 ?���?�V�\;�n�*���G���]K�6!�fpd@O%��Œb���8�\�zn��*��"0����!��uk&���X�=�Y�G�������fK�"Qt�DvB�����(�)��J��
�	���}w��������]Ѽ�?s/Z�K��6���G~njZv=����p��S��˦��V��唥_LѕBy����O}�h�%�B�+����6�h��*wX�\���(U}�܎$(ѼTC�ݙ~
����f՛+�o���6h4'q34���@q�c�|3j8���nGu����̝�be5��M�S�vCF�����)_IZi�H��>��%8��{i�/f�D����:��(��T,�{�%^������z$X�T�'Ђ�[��:���BHK����U��x~w���J$1/�v`���K�Զ#F�*:꽼E���
̛j�4�������W:Ʈq��Ė�\2�u��qI���$�=�aT5t	/�1�'��X�p�;��'��]L�
�r8@�~q� %�N .4���U�Z�U�����W��!�<#2���`�1H�
���h������u��4���I)]�cȞ�wdS�d�|e�A[��E�B�
�5�DӀ9E*,}yt�=��0L��Tn��n�m�2�z�{�w��j��|�J[�O�����IW\�{��̾94�݇cQ��4͈���e/Ld�S�1�qb̷@M`�����,EV��=����))m��,�OV�'A9@S�থ= Af;���<�NC�*���D�OҲ魥�Ȇ3-񩷐��Ut���`$�����ܢ��do���8�y��p���~ƛ��r���ӢRZ%^�@sO�f/ $DFG�$'�g�V���1�BM�4_.I!��-�%���1�&&��S��$:X/�
�Kh*����A1�lڹ�󔠟��W��F#$�l�0����A��;�u/D�q,.����]��$[�?�+�_!p�i�Eی�I�w?;,^�������/�����
��]�6�T(���cKq5؂�7	��w��] 	n����/�e
�bV�Gd�����+D:�@B���.S�����۠���Ʉʟ>1/;�joH��Z<�<vQU�4��t&N��� �voT���ݟ�m9r��Aޏ��+�Xb�K5L�7���	4έ�9�ps	jrvtk�\c~�d�7Ӳe�K}вk�voe�4�a������G�8�_�ʶ��?�����P��bt��vbt�g�Z4��#������%0N�>�~�+�_� "d#�/ГrL�n��4��;�峣�
��u�w)!YH���`�d�����U~�L����.Y����BS?���ְ"�>����ʦ������\�A���fQ>α{�KW��味�~��H46	���k�=�'��:m�X��/l$89��]A��]-��n).'e�8�:�ɽȡ��d���[.�{p���r�>Ѥ7H��,u�۞R��u�Q�Y`��K��k��T����׎�d-���G�E��S#F����cdbkVSJ��a�<Oj�j�$Ng���UlCa�rZ� ��fO�������G��?h�ܴ����i�d�&��Fi�Qf���F����C�b��S5�Y���q�jYaUȇ��!�=�&��i�g4�c�]� W�Z���HS`�t �@��-
�K�ߓ_׬�Rr_��L����r�>G���#�|�S�L�E��G#��ts7���\e+��}?X���~�;������5g����Un��Wne{#>9������$�Y|��v{���~%S���x�OX�˦ײ]Vȩ>��Y*E�1g�ij�hN�����G�F�Y������*MR�{�����Ɣ�>��F4@��!2g?QЍT��x�e�j��M�h�|�(tBҭ17������)�t���!����0�I�p��(����V����y��O8�G������F�o�74���VF��|mtQcT��:/��	`�iK<W�m�j��_vM�}ʋ���p6�My�me�Dt̓�0� �Q��LĳO�KĴ<		i�&q$�v�,ci�6A�������ʟ����}�.b�8��Rp�TR�7��E3 �j�*�߁�!U�=W`&�n��[]8v�vur̰N�=S}���D����8�a-(�M�ݵ�	���T҂tIe7�J��ۉ�хܼ|���剏D��K�����*I2�R�9��@��ŀg�/��*�wSa����B_h�B�q�A�����ő?H�C+$	Sq����`��+n����wi?l���d��Q�l�c#�c��vy���P%-�k><�U�噧��Y��õ>�<u��k�
󉖆v��=j�?N��D��M�%��.iv��v���L���%����^�7s"��3���W	j�Zf��T��L6����xW#H+�)�Q�K��h%�������α��/���'�O.�i�ٲ��~ ���BG~;5BE���l�F�5_�[Cg�O��=��~�ٰ�H��rG1�v0�xU����fK�Ҽst����� 9��K��Y�M}Ҭ�	�W}b'Ƃl�ͅMuܪ=h!W<�F�r|�g.y�����xd��?�f���H�Wv�^\����I���\�78�J,y��S?�_��� l6>��;�4^�|�fE��e��E��@p�
�uU�\c iN{��A.�&_)��ϛ�Lg�e�k�H������ڻɉx�`�輤��!�JC$_e��Cr�;��$�>_N�����=�y �!�ʃ�B!BYr��;��!jD@���W�a@��,ά�Hn���Ret��U���1	�wL�	9�W�	����x�3�.}��|$l��ب۸�*�y1̵ੈ��c�����ޟY�]R���?;Џ~8>�Ue�K�N�@��_Z��	& ٌc.���o�9�����ߟ+�a7��:��Z�	M����^�j$�nɚ�3*��P�Ʈ$�ݳ����9�x�&,���3�~J}$��ƙqT{�6F8�M�v�P�y�]���#����C�fs�.���� ���|98�ۜ�22�ژx�)�7A-ƙ��AJ��N7nv��tِ�����Z?[&����