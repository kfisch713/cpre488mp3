XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Zl��>y�E��K�cMc�����Vlm��dEw�'����G=5��)/��H��n�`�,��[�HoN�m/V��f��<͆�'�pM�#��W}Jـ�}U������EXZ�C���}�}ի�� � Ƶ0.`]\1R�t6l ������	���J��aK����9�� ��߲z�����R�B��ec+P��Z_ ���x��=�X��D��yi��u�� &m��5�E ��2�����"+�����)J
�6v�cIF�u��%��[�{��R�;�ln��IJ����3��2��5�NK�"{�^O���Z޻;�ژ�5����	�H�!�=��d�!�CRAn�D��j�Ⱥ��/{�!X��K�o�K����D=~K��#^\��7�<��-�/��B�탨G���W�19�nJFcO�ٔ_�hóTG4G�@�[�"��s�c�+�-b�{������¿�pS��2�L���� \\�h�Q #@�k@��L���"H�^
9:ŗ5U�������t]-It�z?;��/��k�%K+��O�q"��p�:^I���r1�ʞk,ab���N����3�xP�0.��ǜr%�{sgb
�&s�9��*�\���;��������'qZZ����*{%�e#��=Hm�̿�$a(��и���g�(4�v�O�|���B&'ݵ3��>5&3����R�b[�S���z1���Zh8�� ��|?��@ߩ�(�uY���1�
0�����@�Бr�g����&?����}XlxVHYEB    17b2     880/���O��I�m\�����f	�r�L�i���b\���L��.L1'�i:TCCɞ��Ky��|?I'{J�I����> s�XJK	(gdQO����6 f�Ӳ��
�;�k�䓣�u�n	�A�)�H&<�F��a��^#���m��d�Wl�bJ� �v�� �b,�a�i׻�I���3�%Kk�#iے�e�M�gM�PG�<	Y$����R��ַA;�����.�#yp�0�t��. 8br��&�W����伌&V��E����l#�Q(7eF�����������!��+f�[��m�w�z�Ǧ�2�\5u��'�RP�z7!���+�Nl(.`&V�"�^-\���P*��s�rkW��L��q#���>S#��Z��0��as��O�^Ɯ�2$�@��
��~2a�j��
�T^��ۀHs��s�񐉩iM�:e�Ww�����,D��,��HL��h�����&v�Ifi�%Bǋ�?��K����I�^�t�ؿ����7��Y�;�3����,i�ןu����̪�����N࿮��}Hwn�l���~>т1��1�Xɣ�t� g|�4;A����%%�6>���6�\A�evH�G���\I/�x��1���|�[x^��̟	�B2/���sf�����~�-��u�.�̐�͙]���Y[B̛�;m�u[��92�&����tW�V G�(f2���uEt���c�'��z��k�zT�� r��Hx�T|O��$�c"V�',���/z&�ddn�Z�"d�o�����ʤ������ҵ\(�/D�\��܄�'Xё%�ڏ���U���c?} =�II>7�ɓlZ�݄;��%�Q�y�t�{Ϝ�Z�H�d��~��-'l���I���N�Jy��/�|\!9�os�[%R�����$%A�;{R9����S�OFse�\���B� G��`��G6����;�tE�M>&����;Q�6��!=�R�/���1U��R�����p�8��w�vy{kq��w
�?  J\F��ߤ��-�[9�=K��X���z�V��̤h= ��q咫@z�D�21�i��)���b)��!��6�A�v���1`0�|�JX^\��(�������5�]@�h1y?�I��%���j!�C��w5<5"��٫��uNYf�����s>�,*q��}���!���l-��0_l��z��{@ܟq��4!�pV��]�Q���7�P�4��"H�����DQqP_#s���N��-�u>�0���ush!ř�M�W��JH;bbpol��y_dK"����w�C����+��%'�����9���u׬	u����Q~�����S������\~�h�4�~�gX��G���42%�Zv����=������d��o���5����Fk������بޡ�e�`^��Ž�=<1�J��t[_b����C]=px�%�?��+�D��*�i��98ɤ&����p`hB�̊2X�K �O��P4:l[;�����є�'+���lQq�p`�$>�;Y.!˅�|ŢJ�0�_��M=�,nI����`�8Y���K����@�2��R(S�8h��+�����ɬG-H�ߝBO��cv1�H/��b72%��l�I�6#</��xSQh�����	N=��N&S!��1�����i!�M��k'�wi�X��gh@�\'��Ԗػ�ط�{��@9V[L�m���Z�S�;�Q��p-����	v>�Z՞o I+����.�57�SBBU)�B����3��0�3=�k%bxl��SQ�<����AĮ�bk%��*p�3}X��f��~i)&a�ʒ8���FN4�����:^�φ�t�š�x���һ�\�X�5�߬6���Jx
�Q3;���{"���;W�9F�u]��[��`�D�⌦H�QsX���[��䥘�ݙl�,{_�ޜ�z�.���2��p���������3��!�v�=�	(���'��u��Ũ
�vn��7]�6&H��2/G]ژnQ�����X\��ǅ�7R�S��^��- ��lm:���0�6��@G�(���̉�fFK�f�E��N�	���آ�����G����B��|>�w%����0s�9a�S���