XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���Xu�EZ>�_,�.���q�$���騁�8��)���_n
��S	S?����F;�c�j�'�~:[Y��K�M!l%�t'�����ⲽ�S�5W���Z��:��? Smb�ds9^��|��Ȱ|>�dh�0�:M�1����#��ށ;v�x瀚�D��5�@�Ѝ�f9��Uӝ���Q�
��M��+��Rk��&x�ꝹrrL#�h;������e�'�H֑D�n�1���O{?u驨�����_
�P���3��Gc�M�qj��4�����O3�[�A�S4vg2��ЈI�)����ۼN�۱C�1�o�U��;T�^ͪ ��et�:6YtŻ��E��r4頻1�\1�+��b�2�*K�����̙��v�p����Yy��K^�r�h�yk�%'մ�w,���2������-��\Mm�P���ݣ�%�ڴ����6�z�0������U=/P�Lt\\fNE���#�����80~�;bG/L�Bu�kۯ��U=x��Y�޶ �g��S�
d�E����2d�b��%��<��|6e������h>tgD�ڀN��B���29������mF�[�匱�-���_����P��:}w����w	2�jN��f����RB��=����q:>C�vTR������3���(�֑�3�jF�c��I���u-&1`>U�
�oG���/�\�n��A7a3�(D��Ar���7Q��,(��S���m̈́n����w{XlxVHYEB    2892     bc0h�TcQ�Aĺ�'Ͳ=�
�i�p����N�-�IҶ�g��|L=���1�a����yl�dD��`o,-���N��r�1��?�H)��jM�M�+G0�E�+ZJw<u<Fx<\�O��d�r@08`'Y�oI��5�z�9)&_M[Ŵ3@�����Q3=�ג�/i^��5*�Ճ �z��!��Tpn/�I�ֽv��X��:@���s��T�Ho�d��!q@�
���nM�f���X��@)	�R�A��9��}�S���U�~�����Q�L(o��N��zlc uӰ�ݯ2�4���k�_5%  ���8f�ѩ�8�x�'W�����Aճ}�2���9��_s&���|� ��4Uy`"~R2C�T�BQ�:&��)&/�Z��L��x�<�i誳;�`NQ=��{�ϤZ1L9�U����51�Qfa�L�����<���B�*��V��0V��u�/ G����7E���w����?w��X#E,[4��S�QRՆ;xWiګ���_�s�xe�ץ���%����a����֍����?>�h���X૥,�Z��t2^�~x��K��5�X�I��;��n@�V�n��H�ܽ=_5������];�p{���D���f�bÕ#��.��I��'��vj�^���s"vk;�`�z �d\=�yFB��d�>k!?��T��	�NR�<_��!CB�[תt�J�eE)��r�fRxvo����*�>�re��.�M��8���Va̕8 �7�*�sM�*�5?�����չQ�B��bh���W���>qb="o�b��
89`^8"�8g$yX{����>�"�Xj�
+H�ߩOs��"��	k���L+_�'x���-����0V��5��2���Y�O��x;�OU���$��D�o�'�xG�@��w��4�g�����Xu΄Rߑޒ����(�!��L3-����;\�|mChv��	���M��G(��F�Ft�eY���£�hA �]����y�t���k��2�f��o�����w7;#O�z����r�]n#şՊ�E�SM����JP}[��1Q�� � X�C�'Dt.ۨV6���B݊�I��V0P�4Y]���򙈦�@��/i7�s!�$YH��i	��+ot�Yh�C�`������)�����9���L���+�$�4��G��޺\�~������n��t��9M@�1K߉V��D��-�QI��z�`���_�0�_P�ٓ�/W��d�yܞm{�+��޿&��r0����3�>l�����T�CL�F�J��ǿ�X��A�]�͑�A��8��J/ W���21k�+Hhx�m9�J8R=�jXp������	T����Lڠ�-H[��}��I@��zI���S�ռ��ƍ�>�v�!DAH��Z�.��;^-�GSbGMcV�R1�5�����Т�Wȱz�,�ur��m�}���AV�D6ZkǱ�E��c+Ε'Xɽ����V��g�V<gm�h��Ⱥ򾚡&�O�7�n�@��U�-��)m��06��v!u<�̮��1N������ssD%����}j;m(n/^:�N�턻�r�i:�� �{�<��{m�+'�ɨhzG��=��J��"m�����Q��$Y��ǧ�C��r<�3�$��@5��^��5a�)U�j��}ь�i��a_[�veٵ-+�E	�(��/=�b&��y(M)�jNv~weِS
�}&�=����F�#z���³�V�Ҫי�̼����Ǉ���QP��:Gr=Sp[�,:'^%13\�rz�i�H`�;�T�	 �~:=1HB�@4�0���(���1��v ��Gw��VA	~���M�r9K���(�P�w�����䱣4�������O>�S}���3��J�u+��uv����������كAk96?:�\:_�[<��|⎐v�Q�4��Ȥ����-?l�0��cEk0c( z�19�,N�:��\:�
�^&�r����,p���s��~�ZA~���I"���dz���j�"��C�X����$�<$�V5��d�9��x��Q�T��b���zM������;zda���4������My��=�qK��F�����L&��p4��U<��N9$E�KE�	���J(�����R��o�8��2H�#�ѓ�ŧ	A��f�sE�B�!�ǩ<��Q� V+� ��Ew#��yf�Qk��؅YF���{�z��&���f_� ��)1��;4��U���0Zu����}J�`���v�>p��>L[-ߦ���Kxw�fT�=�0	��}U]Щ}�vQ��@�9K��  �V�YF���Њ����!�s-��A��j�k�[nL=�O��lP�e����΢��:yA��d�]����+aR7�P��BB�aF�
�N�:�J�"�f���J��P^+����?���6��Fe�k��78�?mH�m'w�a��ُ��S�*���������Ed$e���Z��=n�R�5�T�"�p�j�};z����֥���F~t	�Oe/;+��QG؅��oLv5���K�g4~@E��<��qOzDYg���n�V��xv;NK�������)�5�	�����5H^4�d�I�,�ޥ2.ie�(�xG���^�^#��F�%iVȁ�3=|�'v9�&��I���
���2�G��k�@�G��M>?á�0	 /l>(H"��+.��]/�-�n��
a�,��ӥ? ֶ�lg`H��'�`}�!����y�]{1nԼ�T'w�N��W�D㍀��5��Đ*�<g�po��6��dk+��(�RuZ)._���qU�C�3���4�#6�Ƭ�I)%1Qh����d�[U���kO�NXN��7V���i�/E.Cסᥞ߷gD�	_�n�����LO@D��閶��F���Х����m����O��g��rjv��i�7ˌ咦��������8����5��R<