XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���U980�`'��ZvW�ۀG��:b�V��.�eӰ
���A�C�U4VC���O�0Hġ'Y�����Ȑ�Z�R��6LT?>QMh'�a�k��}��+P늅�i�v痘 _���G/�s?�^��
�z0��z,��b1Ϡ��M9v������PV1sW<z:H�qW�"5���ѤG�4�۵��{����?MM}��������K��M��fl�sw�F�-_�WgL��eB�{����1k���Ι &P+�_Bxm��\W��c�E!rC�oBuG�5�j:�ć����G�~=�ca����x:�R���u�C�W���}��4.^}s�����t���|\��V���P6$���<�ߕx���g>���p��} ��{��-\@����[x׭�(� Q+��3��k���/�xv��'$�@;0���Ӿ���a#a�2��ai���QŔ?�@�:�[��U}�Ʊ����%.���e`v�g�#��@̀M~���X�����
;�	�6�S�%�usJ�|�:�i&�����@�`Ӷy��hf� a$�rd�g]X�&��	�m���Xl�b��$/�|�"���Z,���2�[��Y���(�J�W�{[")w�e�R�r
iz(����W��Ƙe�x�h���4Ψ1�tҎ	��C9�B�_@�Z����Z�y��ảO����BitI�1��'|EY���)���7872�H��+Tp�Ӥ�2}�Z������4�t�يAMe���m�ֱwXlxVHYEB    5fea    1830@�^'Ɉ؀��-��
����R<�x/�FX��>�R`d؈d�M+"o(�P�H%�ך�A��xP�D�t!P��P���� ���ˤ����`b�\a}�y{y��k��L��
��a4<&osV�nL���
��U0ŧV��nR�a�`{�nj�أ��h�d����m��@\k0�����D m����pڅ�NQ�j9kA߭�:��qdJ%�m�8�82���y@r{��E�n����d� �6������.L8{ֶN;k<���j�Q> G=m��=��I��d�d��i�Ps��!M���՜>f��϶Etl3L�����m}5��D�R%vt��JF�N�ۍ���VR�`��@��uT�ºU��&� T
�E�!'\a����F�:���+�bi�ة�K̞LV�=Ө�?S+�3v��xn>ae��)�����c�/�U�����#>��U%���%��TI�E�ԔP#���ːmj��L(��m�A5�������������������m5����ny9����k?��`m�Z� ���'���WH�/�W<���~o��R;���I|Y�0R�lK%�Y���C�3��U�c��Z���>��U='^8�P_���*��{d��-A�q��ki�
��̛�}%�R8H&���.Oae(�Z ^[h�1<;�{$֭��/"�SQ���?�2�f���"OI�>tð��L�TI|ܮ�Q�427N"��䒕G��mA�n2�Tr�f��*�!�[��e���9-�+:Ɣ��Q�xl	cb� �|�v�k�b�!�3F�(+�l��
�E���-�"�F��&F¡<���� k��qݡ������}9�C���d��*'r��8��E�rf'��;o�'�����:Ь
ܣF�\��tܹ%�e:�8�E��}�srj��=	Zu���l���Y����C�m���cf'$�cX�S̊x�Z�]h~"͇خ\�<M�ӌw��b�P�g?NM*��2l������s�Y&���f�� ��G-�
�Ap^�.����yWY b=E�V
Y0�^��� :t���?t�|2��g��}:4���90WQ��~o�͝mGI�;$>?i2��ϛ2=q��Ҙݣ����,vZc�M��~"X�?��z�u���:L_���QX��&С�1�ڋ�𵃉
X��%�\��@)���5�7�?��+�2nr�7�c9tCN+#�KL_(�v���~���OF?	�ʳY�ј��.}�1Zi�]q�Zk�c�#HM�k��I�0B�v*6����R�t	i���Զ�s�]��C7&���g���Fw٬�`��0m-/�JC����l�x`�����V��[��g���4Hx�/��_w�L'
)n��"�5��fg�`I��H˒KS�5�"�"�wn�XC�ʢD�f^�>�T�`��&삼���?�[��D�4wl3p�ʫ��@b2AY:1��/*�E+��DZ�&��&���B�w���b9.\i�==p܆n���D�h�Uj?{����A��j���
��W}���-�����Y�Ia�|�z��ޜ���e_|Q�ik>a���%.��۫���77��+@��1�Fҩ/p@�r}�1`�Ǧ1�9&q��Mglm���펲]����|�p���	R�).x�.?!�Jm,�"�Y�|�nM����-зV��>\�uր��t��Z�.�ߣ	&E�BH�ˣd�Kxv��0��˯L�#�9���66�'o����#^�)O�s4�ձ0	<�O��8�܈�G�y&�#�&�!L��7�ː����d�߬?[�%�p�@LE�yĻ��c�bQk9���R�ė_Y���6|�Mp�-1�0)�k�|z6���BI* u
7�Io܂| ���?W�oǬ�2a�9B^-s�p~9_ŗh��p�w��-!5�Lr���>�ț�^Ϥ.�@u������#�qN�Q�M?ʔ���m2������@�]��fL�#[�,�q�J�f�V������0�|���Vh�>�d 	�ʍz��}��|p$t;פF��k��_�����)����2V�3���+7� �Y�zo�����2��a�u�*��j��v��(7dQ���{�m�>
`��&�*����]�4wUKE:H^ԛ�d8N4�r����\���ƶ[CC�B�:5��աr�L$?�E�&w��לGݍz�w���C����nk�ZA����i#;���b�w�#¢U�"�vR;�Q��Fa���N�=�bm�i��Or���_�a*A��C\G���<S|ŗ�%q-�IRNh��Ϧ|��;{��v�U��T�?���P��@�^�!&�v��E��$'��s��akY+������Y�#IgU9�|e�j��0}j�?�={��Xx:y�2����2�J u��%U`��$��նsz:��1+[;B�Lo�k�+މ�Î� U���s��6�y����\�n%$t��wZoP}���l�#%���^[��-�.�I;�	��R��9����^��.\2�b�,�0�[A D6-��JN��P`]H����G9�k�4ԙE�G�	��Y~�(�R�ÎL)Wy= �-��]��&�k��ɼ+5�"ɰ%lWN��rj6g��"��{ϞC��1�^�D
M�ZŢB쒋'�+���'`�6d�|��s�S�D������hH1N�/.�9"N�Uh0�W�v�^����6�`E6�=�TV�Uȿ����j�`<Đ�6>��{�2����sg���3b��y�|n<z�~ڊ[y���{$&��<��b4q[|��~���멨�7��ab�M�.�3�S�R���Y��<�0�R�H�4�����-�18��L�~ ���g�"�s��p�\�Q�\��:e���/��G����2�H�~����|�bc]
�_�8��?V���< �bɉ )�#F呤cGy�$GdC�0���qq�¸����N�mn�T�f��l��a�`'V�~^�ġ?z��^w*1���hxއ���]������7���%�i�iZW���ô����f�Y�曢6����w��Y�x*H�&3�-~6�W3%f�4�4�{ڔ���5MH�����=ʜ;á�:�*Or[]r�7:�ع�mkv;��a����g%B���W!�y��WX�8���kZ4s���=0�NU;�����ފd
@��������nD�g�W<Z�����au�ޖ��	�(`:@=���}�M�߹�Y	b������%�Ͼ���ӷ�'�iz��'�J�5�}B'��8�H���Cy4�	$���^ �\6B����6�2]�?^�΂!/r0l
FC��܁��U�,�S,ጣ��T�+nY�YR+}Z�'�����!�c؞�&ea���=O1p�K�*i��A��`�q�'S��HK:����Ν�Lcq��?�)쓍b�F���١M)��I��K�:�/[RdV�ցm]I�oXe1HE�h�o�Dn��˧[n��[e)��G�JؒP��98�h�{gڙg�-]����Ő?���y� wdi���3$KQD��Qr���FH���i����=use�{8YìS�_���ՠ����pw�P�W���^��<#O�<Nq�c͸ �ƿ��$#7*�śp3G.�i�'`� u~Q��\_)��'9/���CE>�a;��O/�g�f�y�4DK'���U�k��1!\����b+^��~��̑Z4E�#������9�1�v�$��Lʹ�5�v?�qsd�\|9<�������5�s��[�4�g�[z��D󔋁���_�_>)�ф�7&�7K*2��.��D�I|M���B�V/����YmH�N	��ޢM(�E
݂Sdo��s+Mv�adm+�ݩ��F,��ܷvUo4Fk@��g�F��?	p�;��}m�'�>¬���?���:��LBSh�ZI�t{���	\֣m�]��V����� �)>���Y�>����}Im���y{��m�,8{����H���UK��aB+z��G.|W��fS�H��c��xQ�@�T�G�ҴW�jn3���9��}2A9��x���ڶZ���t����lQy�2W��"oB���o�mn��Ix�O]*G/���f��u�q��<����&�qp���-9��8�ʌ���M+O[����'���v�aұ��D%U�PW�l���:$ܐ㰊/R�<�p�s�'.��v�h�r(TO�X�D&��7"��w$�t�Quu�������v��G��S;�A��:�˲o=1�qv ��ޛ�E�?ʧg���+��.P�ՕkE ��^	�#&1_�_I�$l��?�1z(GǴ~W�a��"�媶��sg�-rY:6�7RkR�P���9;��No�3��/B��q��]��'X>�\1 L�6���f=P��U9��(-�^O*tt���Ƶ%ʨB(G�m-O�+~�J �v�M�E!��d��_�Z���0G�}=[�pyˎ�`�߀���g�]�`$��㎻�<hė��s4�<��� 
��<���?5�S�F�/Pԁ��P�R��]ߴ�hIu�3X)%�Z3�='�`��5�z�0Vp*I&�sK�%��a�u;R�P���vg6�cLv�[�9�#��.x�9=lc!�����t��S$刟UZ�`ڥ,1e.���i��	v��[�z���S8VJ��q�aퟻ|����O^r���7;	!B�O��8&��\M�rL���Y�%8�/�	�=��h�s)y�?'۩�6Ym$�OwOf)�JYWO� �Į��Z4��~$A]�>c&�ѡX�K�)�s H��MGf�Y�����S�_�t	6bf��:i�υH!Ɍ�Y㻻���lI�T_$fH�Q4�,��/��Lp��E�nR_6�Fv o�$�JuSB�1����L ?�Tv���x����JF����p``P��,b4������
�>��BaG1�!���<�e�Q�`w1�|�"ZN>�֏f4���ꊔ�?P6+Wm��f)���S�zA�Q�)��:N��S��C�;
�8�*�H��7b�N��3
��	� Ќ�#=aU�Zq�7��&^�9����A"����BC���$?�!��;ȸg��������<�t��2��ɋ�A?��S�5�= ��,;�&C�c�S�3��)�4Q�<Q�|Y�+x��&���%�s7���]���ѭY�
1IT6��[eҎѦDu�黑jS�7��w'��,�Ô�7�%��H$"�r�S�Re�+AҀ9��g:�A�i~�ɰ�M��:�~����������'�����Q�<^$Yݢ*�9G�KR�P]t�ԑr�j� ;aԭ2�x�H������U������jj��ZIמ� ��/�H|� �����Y��Խ��Ð�%�=���*2�#�¿~`���u�{�v����r�H���NY�͋A�H
��h�4�Fx	4�s�4��Kg~z&*���w?+KN3ǔ�%o4�T�?��~�5�F�s�t��
��X��>@��d�J�I	sL��a2>ٱE�3�[T8 �xIu���ؐz�z���s�\h�Q&sK�ު9�c�I�����ڸ�.*���2�ՠ�n�����r��'�h�������"G9YȠ
����G4�վG-$k���Ȍ�������c���x�CtY+ys�b>7��T�R>b��/���n�8��>c4��Z�<}@U�������ʬ愤S�%d�����R�ߖ&0{*�G��-�/�ׇ����~�9PFL�����)C��w��D�GD�΃V��T:�)�KQ��
T�7LB�`���¥4�	>��w�='7 ��(��6t�e^
�;H+H���rr#���
��R��"nF=�����Ah�����s���*v�i�@�q�߁��k��\��	�`��U<G}���.�LŔ�{`'۹A��(�ǍZ+0��t�Į[��eo���!�:���9!|Q�����,�ue�f��c���xI�x���@X������J��a�ŀ��<:(��A�g��拉�T���LX���̪���|U�3JJj��.�����J45� &�ܞ%��;j�w�q��g�C���Wm��������`m���M*IN4.�H�N�9�