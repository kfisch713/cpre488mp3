XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��1����9�hί�ĩ�o�[��-��$���9j�6�)
�xj0�Zt�L���]|��j۫��⨆��L̠n#��ʠ`x� �^��ED���rS����r ���E�J ˽���2�2U)���)jdV,#�Q�K�"m��]��!��~;�p@6@��ŝ8��q�������NWd���雂���gib��@�O����Q����	��7�����y+I��)>�#��雭:��ÿ~R�+��������X��[��>�\n�S��3�yyW�Gv)7���UJ{	������cA�3>��l�L����C��v��v&x%������xG0����w[��C�u�Q^��a�j����/PQ×�Ek�B���k<IP�"eǀT����+	B���f��i�g�k#�\�1�d�K�V���[л�ٟ%���P�G��:��'�8�)��}��0�(�i�(�3�߾�Dq�_
�#R�t�3W��e:C�H��QQG��v\��l��E�l�J!� ��KSp�\��կ�r�$��>�1"+��ʊ�T�걟-~�|��6§��:]|J�@k�|��
��|i8�� %�^E�5�V�T���9a�'t�,���@\I�uYB4Y������[�Tl��i���!�ѕhV���ĂX�Z.�$��-^|�ߙ1�>��{]�u���Pf�"���?�z�l��l�qY޴�Zh-��2��W�|��
;-�k��9���aF�p��;�t��!׬�Q<�s���±-���m�XlxVHYEB    1ea4     920Lz7e����"���qC� d��0uy������^����1|�0$��z�D�j�lhh��CS�B׭��E�y�/LN�;;�	WM@}7�Cj��qx�P6}�N�e ���]���7LY[bV��9D�( �$��I�`\�V��(�L��L�,}䥿E���z#�5�Y�H�x,�y�Ϥ|b�qȝ�(�cF��L��8����W�3��Q�wx��o��������t��6C�L4���"��LU�|w�J��R��3����������936�\-v�`��z�ES���h�$�g����+/8y2�Vާ�Ւ,�6C>Ck�óx�9aDd�̿l�x�JAf� �KΛ>BrO�%�� �iX�U�	��JZ�9{Dɞ��C�b���P�
�[�}����־���^&V�[r�4��8����2�_��n*t�,�j>/!�v�;.p幸F��x%�ʎ��m���DU��wy>+HI���1tEL�(@x. ���Y���S��R�b���"�(�@�|�\Cξ��qf�{�����l��د�RO��	<�e���%#�y[��%T��K���<��-@藬(���W#�*��wKw�m����=kF���ʀ��~���V��R��ć� J!�����t��%�b2�VowW�k�L��B��<@��=WX==��M|�Y���D c�{9c��#|{�,���l0�e-¨��R�WM+Q[�Ǩ�����g��O���"*�Q�e��F��"$�!�R�ҥmL���Z�3�3��
���Tt��L���A<n��&H�%D�-�wRW�zG�����{��B�$���3�.�Fs���ɥ Y�����(�^sO�z��<a������`�u��YF��&k��b��S�[[Ў�-�"x���'P���Q��%�Ѱ��=ĮWm)��{��d���R�i�T��I����f�T�k���{e��	�W���/�
�6�F��h�2�!��@�g$Go�+�;�K_C������1��Q9�;�u�qz'�B���j��*������mT�ԶN��*N<e�s��zK�� w��m�-�N��GL����/ϣ��8��������]샹=��_&��l_�v�)�]�M��0�h�_έW���a�a[�L�=�l�@�$���;�y�Pk|/���ٕP�����IzӜ�Cq�+��K�T׍��x�)��/A*�+B6�#���>M���E��q�Ml~O;M
��Y�Y�����ŝ~���I��dN��ϯ��D��=�Z����fHe�� 
�j�e�xmPHbfz�xo������V�ǽ"�	�2�~0�HE5P�_���	�U�1k�\L"����@'�R��c�tJ`��d�*Y2��q��!5��j����͈8��q���?;��*���mg�}��9���B+6_��=�0y��?���,�/O%m��`5��J���,��z�l�VX@�=n3h;6cS�L����j����!:>�.X�[l7+������k��7���3�gӏ�� "�f}�c'�S)�h��T������82b ��q{�����λT��ӿPN˧r�&��٨��4�'xAP�h�&u��yr�'�S��A�C��)��ܼ�$��E�[vM9��eDH�֞�t6���
�:���1&��+���
O^N>$���ܛ�sx��"�t�&)��/�{��
�L����+���y�.��ϧ9��o��J���b7�/�{Ni�Y�}We�q��獴J�`��*�X7J�ó.;\T�,r�ѭ[Ȯ�b �-�s����,vī�om���|>�{g�\K�u�����Y��k���$��c�c�\y�J���7L,6طZ`Y�HN��]����32!�,?܋���s��g9����r�-�:�|����Q�d2m)����?��t 8����f�`��Y�$�^���[ݺ8hv��7�(�W�z���x���@2�5I�e���sz��+%r`/R����:u��:̔}���C�,h+�-?������%��X�2�����ݰa�u�p�hA��j��K�Η����a�?�tփ	@�
i���e�Gp�,����r8+fV��f�ψ�����5B�O�)�e�=�� �K;�}��X��β��(7$W{0�?/0�L��'u���79́la�,����Ǣ�(Hf����� Z�W͎�qɂ�n�W�ʵ�7_]��NY�	ĹM��e~kZ̉Q�8��9����j���I���MY��צ��*�d.nn�<*&����gC�ϴ�HY��*>�s�ahcv�G��^��