XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���cQ�8�Z�/��iD�35�sE��nA���������'@�k�Y��.�tio��N��u����tا���*d��abլB�0�-[��î�tg��8AOR=�%Rj����v	T��3�Ҫk���j��!�]j"�aڿ���rֹkm�"r�����i[3����vЋj�]-����F�k��J��k��M����a+F�LtD���=��(nG���^���`_��C�̴!�*Pjj�M���.�'���K״j'�X�=�s��NT�X�X[FX�j-�>��Qy���~�1�)�/�&���Ώ|$���7 v�a �Yz�3���0%X'1B��u{��-r�׌�cJ;��[�c�~�3k�e�O ��v����0�H�䛍���P��w�p�}tcV`�<�,�B�p[����7��;aò�-���y��@"Ν�@����'�\��H�E�HZ �x��$�C�-F�Z������@�:���w5��Yt�n�Kd �5��]�y��O܈�I{��b+i~��;�_����O�bP��$�8.8�b��E(M-��lg�S�y�M�:��$�K��W���0,LCbԓ��!D�\�;ޛY#�RFƚ_1X�}�(G�͔Gv�t�	]�����Mo�����S�w���%J7����K� ���Q��#Mޢ�NMa�1:��8J����қ	=��
]pU}�Pk�@�6��ݒ5�[�M`�a����θf��tq�WJL�����XlxVHYEB    3b09     f80���@O�#.1��jln@�r��_̫��:�� �M��� :u�RH���5!�1Ku��Mt����I�X\����?�ֶ�d$��E�W�;���Ү\�V����R�=�<+���)�d��>z����Y)ԏDv�2d�˗@,��'�5�=��_�ua]$n�� y7���1�ِ_�?�u� 8�"��1ߴ� �k>�57A�8���T�'��Bba����|��*U�s�a�=���L���6����)X�Bn���>k�ek�O����'m���P�)���S[Y$}��vLͽ��]t�Ů':��C��I��J�G��j�B8� �$?�d0A���g�/������+�'`�~�1�vjR������lԙ/����Jo�?[dL#�W܉��n�qS�J����h9
�k�H�M�ٗ��uxrjޜw=�	nĈ`]�B z�E�3F�����Mwbg���PBDm�j�#����]B��䑪��O+���N�4�P�o���ђ�LNT����Vi	'�3�)ܤf&��_������*�>�+�JM�V���{c`�O��@�hF������G(H"o*�Dӈ�LT��K?
2*��濄=�<r��[h&'5!�J�]�.�1v�0��y�i�=���"7�8c1BX��X!.��Z��5_VK�=V[ˑ1�]!ϻR��L���T�6�!�h��0�x�r�?q�[5��ooa՞ɩ�[� �֙QlP�6���{H�ק�ק\�x�
���f��h�_P�(�u8���)��_�����Ű����4�nv�{�y���R+�$���]^�ʳ���)�n2��ߴ@�#���V�Z"�>�K��$+���Ӵt�9<8�/��T7���{�H���+��艡g�3��P�A��s�`6|���id��(1F!s�]�r�\��n�h$�6KO��k�8�M8��Κ��ع�o�ʎ8m9�#�U{ ��$c^"g{�������!#�^��R�Rr���X����� N>��'�T�_(ma�$� ���xU5d��Wv����FN������P=�`޾M����4�@��(�q�+����
��L�
J�q�j����	��E�[NG�L$����Ń�:�}N��B�Q���Qj��|���gDM� c�?��gڽ��,0���ͼ�H�����1�Q㊤�i<'o=?T��y����A{���&�
���F���|e�흻��Z�.�x��:s��ҋ�e�2R���'�p+��_F���g��x�M����Sb#%��AHe���b��3|K��D�醜9��s#��}n�,g�J4`c���^�S�dA�(W$�zK��o2$��f�����	�,\���"�ӑ,g��/�GolRK�>�w�)��0wQ9�Z@A��%&o�j���O��g���@y6a�M�Y]����?��������2$�>��&��B�(���uC��@ǳKBʭ����BWL��	��lV���k&�����F��������U�8!��ќ�I�Eo����<E��8zȖ*�8i	���<��c�z���i�j-�-��&7�p���� �a8�7<C�W,B�m~F��p�.�b���,N1���j���a=,�Zzd�En��~�`W�w�G�m��,�p��&V���b���r��YA�O��[��K�+|�A3����6*�d�����#�B��T��Ԋ\j����]#Z2���m�ر�)m~��9��>;t�,�Ml�S�,��-�hA�'H>yL�p�T!��S �B�6���?ȥ��L=��.�.�e��4�7Y��F�To��;:��d��V��}�
��g�1��.���{}��Q���Z��1��Л�@�X
3Q�����4m��A�y���/�_X�R��(n���_�;h���Q	�!M=UK⒙�/�JU�?x�Ws�m~��9әH���k�w�����w.��5�7��c�R!�w�~G�(��J�{;���|~IN�q���b����B��~�T9Nu�J.h�[�C�)�`���gN��o������^|�/B���n�3������|$�=���3�
H�7hߚ�K�Na�{g<CcoBXQȯb{��H�"��[6%kHȢ�*tˈ�A�?u�NxPܧ9�� �c�o}}�Y�S����Ͷ������=�����);�oX�M�4!Ow�O�����tX�kg���O����gf�6��U�^K9�LS'��	���ђa-9��L���Sa�%d�WOL���p韺��4��9�I9�/����i�Y \�)�Ue��S�$��Ȼ���|~�X�҆�Q���n�ize�bS�*��Ĵ3{G/�f�D!��aɟϠ*�Ԁ�U[�y��j�$��-��T����0��Y`UB���5@h�	;i_M��b顡��1���������f^�"�3�շ�/�o%(Q2�#��ȝ�7-4����_QP���r.������>ߥ&~%-��"`Jk�Č�vꪣ�T�ϫ%�W����`Sz��c��6��i2?�Χb!�AT�J���On��a ~����i��{��b��3�w)H$���)d�ax�u�ki�β2Ӛ���3�-V3VaWbj�!�|*r�r�T:�&y��r3�ׅP)���YKF�g���v�o��7x�a�ʲ2�Ww��Z�q�źk&?)0��6ӶELn�1��'oCo݄��l�4�	�C$b��EE9��S��z��yl2��T���S�i�\4j��o1W��M\_zUfK��t�C�ߒ�u�m��kN����I�'����M���u���X��ȡ�������.m���J`i=D���Ϻ���h2��`�
=��i̟�\&P��\t�7EN-�>_w���+�Ox� a*'y�(]{ѩ/�r;�UA���9!�-f>�<��}?�˫��A�&�g�Wl��)yp����'�e1�l�A�VHk��Rj��6�Ɂ�Vp<1�
T��#Q����=�g\���V�ޤ
�����Lt��Tp���'���є*]��|��䝛R̡B���45D������p�^��٪5c��ݩ!����g?u*Bݛ���u�*��R[��L�Q;ЯMJ�,�)i�$s?k�5u���S�y��{����`�dH���������6�bV(~-�7^v�%�Ȣ1c�d���4������X�fT,����|�L!��բ�i����a�L�V�4��Jѱ�~dsH�j�0�����y�9�O��m^CN��RI�i
1)Qf���Dg5^7���ᝮi�|A��~!%�'ێIƩcz�o�$#�z����t�	���S��G���V=�=vD�:�)��"7C������� W|_(�z6�@���j�.�v���L� �ʋ�F�(�Dv8�zG��c$ydD��̉k������5:X7�Br_�\��� V#��F����V���������hi�і+�������w,!a F�9mh�~e�J���Ɩ�ٺ�1���c�O�}�n��:�o���)��.�u샑�{?}&���K�~�ĂO'�QO�"�(
{����m�?iu�������M�y�X.��/��7�^��17ݞ��g�|sr�K{U�l�M�X�2&f�B}�I`1�$I�E�tN���j�ҵ]��[F�������4���l����aE}i/�$�i��7x�??0�ʇ�}+'���:>1��3|(��kϑd��~/ڐ�\D��Q`y	�N�T��\�}�z)O �g�������Aޖ$�4vIpN�#F�.$(�7���re}�;�#���[�F��Y��	Hts�jx��b]�!X$�p7���ӝ��8�.��NzNn��,��t
&�Z�9�`L��o3ٜ��q�Z�j��7eɽ+���]��