XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��I� �H����-���К����	��-�i��2�sh�x����Ka��a�?�b�N����RTK��癢���i�N�OK����u�	��A�YZY렣�u�'�O)����;F�k2r��D�n���&5y����r�F����;{ "
]ڍE�S;�ş�$���vM�,�N f�"���;�E||^�^l�:A*VyP��H]�P��2����#� �;��.�g�Yi��U��ح㯃�;�D�A�"���Q�p}�e�[�C����y��l�q��l&|ۢ?/	�Լ�=�y�|a�oG��h�r�D&��=j�NpG��~W:r�K��p�̟��0��I��A�,��z�������]��U"ȗ�u�b��<�c؄��bp�ݭ^�"4�����dOS�����:�G���Ol7���H�s��Qj�	�6�?GRѲ����k+[Z�a�M~�]Z��~}��Ӳ��7̽	�����Ľ/ڄ�r�h�o@8����O�
+�ʬ��P�d^,3[J٢��#�a����og�+DL����?��21��_�����R!�4�/c9H����3xN�i!A��n��X�s�y	�`�݁8����}`ӑD�?�rއ�"�:[��b1��42�8�aB��`���.���fj2���������*.��-�Yv���xsA�j,��س��S��[����y������zC~��x�hl ���5���i� @y��� ��ȼ�8��F����#E�jfEXlxVHYEB    7265    1660�7Ex�nX��8)V�����*�/����?!�~i˛L3���#	�*����J&�i�jJ��D�%Vԅ�d&0�(��DQ��&։M�D(��WdONb_}���`�jH[
d]TN��ѧ�fq$����	�o'���^͒���$x�ӧ8�^�����$�ΌK�l�����c����T|�1ƪ4�W Kt�+��a������:�K�(g�B%;��/_���	{�*��J-®��s��������Z�I~�����n���]��YɆD���^8��;}��R��~��ځ�;��KζK�������+��\�巼ې�`�K�j�8
DS���!P��ԥ0"IԫX��`ţ��S<|5od��=�H�cO 2���*�S!����\�N&apM��AX^|��
7����D(紃Ỉ~}Ŝ�
BܺZ��f&�þR_�B�v)�G	$�N�xǋ6�۬�7���klwa"�rr�����CD����kZ>��q�&�����$�-�pr����ƩrUoN)��tA�M���MG��)hb����HMV�Ax���1]��u0�����n� ��à���X]�T�^��cC���.��3�*'���7	��
,�'��{!�F��K�3 ��"8	>�W�lt<9�S'F��QG8���e��U�1UF8AF�PYƅ�)���<�U��"U43��3/��B�I��������J�{�j��=��f?�=�E���aMC�6ZmS~ b&�4���s�.,Ba\�� PS+�nt��)C��	掿�(kC%a�yZd�}��=Se��ζ�́\1g��wG�
j	�C���z� ��Śk�)B��?=��h�=�5wR�S��Ҏ!Qwd\"x��%�=��1,�Q�=��sM�^P4���=���]�����m��t����(������/A�~���Iy(���D$q6�P�M���`�Y���e�@��s�>��B��,K����qw�?�x\��KtX���ˑ������USnp8��f�8��ǧ�8�G4|�k�!*M=,4{�R�ޞ��)�3������[��^i���7q�L'��M�����I�Z�Cc��6~Wk���Q[�Y�_�a�����ȇP��cca��D���<c�$a˒%o\�ͨ~�7?'���o�\�w�������H��Ǥ���XN[�����F��G, 7�����a�H�Jz#�[  M.�b5S5(Ce!Af��o�H�(W=�2��i$f�)H؞�)�A���=1`�*���|�W�:�q8��,1�Ke3/�Ǩ�$��O��'��D���C��:��!e���O!�>�4҅�7E2�h^.�gs�z��pu�|���cg3��{��$��af��|)�el EEݭ��ҙ�ὣ�"9�z�8��������eͱ?g)Ġ�cT�S.�M)����m@|fq�Gw ����G�FM�wL��9/�e�1�ݤ��m�2ꝅ�r�3��/���K�c�B$:,�X�����@�pN��}�[=y������?��O.p��vn!YW��=\vu$I�@q|�[������ꯋ��F.y��r��t�,K���#n�;�&��-�F9�p�8W`�I;T�0	��am��İ���Udap�uS99܁`uد�;J�_"�@��LtӺ_C��K�Y�����
*�k�$A���ЃҊ0��؉/x��z�B/�����V,�rK}��x� }��
�>��1w5`>�5;|[��)��溑��Cs���6,�r������`&��U�*XD��&��?JH�e疌����ƙA1^��~8��xwC�B���Rv8����)�\�Z��A\}�7���*Iz�E���̱�����;�|�H���^��M� E[��q@�B�6֪v�&�@<������f��N0��,���?`�cW����="r����'�Hҵ#����Њ����aW��1�~Br|N��I�B��cC��`S�eR�S��%ӌ���~j��]Nv���╄�f>��-��&h����s�a�g
snx��F����"u��9���_��kH �N���3�b��+�����WH��͡�-!t��Q10��M7�{,����l��v�F��8�7�0��.5�+]�'J2#![��a`�ϖb����,vb�[Y8���Z�� ��F�Zj�jI���V�x�q?�I:�c���KvZ~��Zo#ф/���=�y��T��.FD���y*ܭ�+fJXa6Yk�%
��Q�����u˽ךɈ��`��<n.����Gv��4���m��e6���,�LM��bP�;�8��tq#b2��*���ҷ��@�}���H=ϴ��� �VN]AZo����=���/#�ɾr�c�Ice7b�P*�%tAۙ����B��UG�7�Kyv�4�18EnJ ����O�찭�\��w�.��n�0��1)��mM���V{�����/A`Z+?��Q@WR�!��-+��l���#/(~�����0�c��rF$�ʌ���IHJ���]Ei�u�!5�H%��Wg(	�~S�({�u#zlDw�-,G�G{}��=C�@.:�L`j���*�L�5�_1~o�J�����<Ě�ްgl��Q��82�<��M��ҩg .7�� T��u5���:%�|�:�H���Xy�h�U%�RA�rQ�ڼ>��9�Ǡ�ws� 3
�say�>�f�nz�.a����buBu�t�v��(�Q�K=��*����M�J��{��?"����Rؠ�	�^���Y`��m/���:yl^9hx�jڠ� �����8<�:��1r^��b�C�p��G[��Ti5���f���5��-�0�2�u�Z��O}��S�&�_��8˱�%&z^���f�� ���ז����?�8�B/�r����z-�;m�@����O|-C���O��S�>���lO���v="e^�'?�;��ٳj�Λ�E�8��/6 {j%�GT�h�q��4���5Z�;$�-�߮̌2���yu�F��M?���/W���Z��|�g8���rLِ�#34��(�_���I�*SD��q���"�t:�O;F�jT�b�^���E����|J$7�����RHG���.�{kpp47��4n���`=�QV�=\�c0�ҡkӅC�y������(�`�M�� X}�i��1��(q��~��	��]LڑU�uM�b���"'T<y7^˿{ײU�D(&�j�	~FYC����,���M�}��G��'pl��7E�����N�cV��"�+�U2D�]x����G���v��[V�V�ʑB* Z�:(����`�
�н��GtIע�>��Rld;��A�5`�A!*+��B�%�h9y�R�t E'��U�����(�f��2ھ��@���K��Yti�	Y�m��v-��b�v\pm%���J0�S�����*�����`��}z~^͔8:_z��� ���5]T	{�"���������'����'�d���M�o�^B��A��V�F�7ɘ����PQ�(����6��z�C�Q�(^��Z<5O$�"l�oh�S]��L`�'	]qC�Y������9����W_*�36���j��8e��Y\4��hn02��
��4zX�����f��U$�!������j'.Z����d"�ܒ�F��9v��GVokKJ���S՟ !�hB�8�퓹�f��T545|��W�p8�=�nHH1슕�SK*#ڶo�"��tc��m��:J���H!���
���y��|)bk$'�6��<��nh��Y��sDZ5��|h�>�M��jl�i~���V�����L�%�+�Y_�T6�n)�4�%2�h��@o;���}ڏmQ[��N��hGNr��\*q�}�MԷ��<6�m�!�f9}��L�e�v�޿M���u}-:2�<�9.�y�ΓS�ǡudp1�ΐ����ǃ�\-��J(��o�f(��rT�"�����])�iH�a��7��2"|2s9���F�p��GM�V��
�W�-^�PCC�Y��%�=�l܉ s`�=��	��-د��
7:��e���G�H��)dmw ӏa�Ӣ]E鼿A-���ם��|�p�q��f[�=�8�i{��!�K��X��`���l�~Ώ�*B(o!	�Q֒�ĺ��8yxy�ӰB�I��F�V�P����*
W����f���%�\��h�VdC-�gt���N��{V���[�Fϳ/ޑ'�A��t�h�)!IZU4���Ψ؟uގ��yW4'�VOɻ��W�h�2���<��q�S�]|�uU���_~Ggx�L�R������/����.mȱ�6-�+�u�x*��9�X;aCM�	K���^xg���ȿ,q�,ԙ����Pg������6Y�y�޾*�Ʒ+�qy��j"zy��F{�A͕b>v��wV�Dw�=�9�Q|�L��D�hn]�YY��Wߖ�)[w�#8�۞U^e�b���d�_��|ڦx	S�5*����u=�M=��a��@�0��(w2���ÔVw���F�U�'�a�s�m��U=y�����<�����������Odb����(��<�0f1چ�EyRU�?��%O)5��>M�$���>�Q�˻�<�3�j:N#Iwk�`��h��y&h�y�������#z�_��f0z7�nex!Ù�L���᫵�P��;S�9u�8��I�K_��C(r\t��/J��{�j�lwd �IH�5��l:d�@-Ph���uW;��5�ο9,���hu�'*�7N�7��ۈڙ��^k~�H�kv6�W�y؍� Nc��D���]P��"e���|�8��n
���'�:^��T6iW�߸��JE�̓�S�)5��� �謯��{���Z�\���N����oOJ�������p���j�1���Fӧ�v�(�X�����󍜉\z����'`���/n��3�y{�.=��nDUo8^Э�yEYÊ���'�[P�� ���T����Q������~PMp
��x�Z�zC�Y��I�1b�b�����P�4�(9���1ll��D����a 2k��=:�ac`�K��p���Y1��2��mm"�9��/�=��aR�P�*&�wx�[8��i����{.֭�%���o74�9[ӾZ�u^�w���:����v&�t�j��.���H�?�	Z���W�T�n�w�q��~�b݇�&�?��/,&Onp�*8��Ω������`<(%�բ�~��b<����s�	'��k&%J>�Մ;��2d�xg�B��_x�7k�����0�� ��V��\�yff�n8a�%L�-<��\�R1&�~�iD�6�
�c�y���������_���߾�77$��T]AI��P~���;H�y����Ԉe��o�8��U�&�����~7v�=wu�5w_)�cR�n)t�+��8ށ�A��^VqT��N����/��L��4�'39{�r'��k��v����
��
�.������(Ԥ���t�h�'�߯���8��W�z���\����{1�2�Ty�]�樣�VS��V�P��0Y��ݎU`��?Ih5sƓq���u�^���*��y+��-1Μ�ZC�`L�p�]��?A,,���Z�$����ؾ�r�7���=B-����