XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��q�r�s`��CSF�#��X!�
/��_�s;k2#vS7��ww�=�/�J�h6�崯G�T��8�<��%u�;~>}�GD��8y9&N���)�^W�>�=x"����U�ߖ�,��^��ǦyD��t}*�M�d"E"��}�f�%N߉�v
��;BХI��h�!t�tvR��ֈ�<�-��CW��ԕS�������P���|�g�|�]:3~�t�ye���<��tL��wdB�X������ѵTT���5`�OD]"x|��u|��}H�I�'�s5�9"��n��B����7�@M͈�c�uZ�Ŝ�}�r����1>�6\��#�{���{�j��]�A�)p���&x�\-����&��A��	L2aaa���D���r��*�G&�gM�fpi�u��#{B6��/����%kY�M9`��e��,�I,�s�ʛ�ܤ?�R>l�x�rU�lӵQ�l!}����2ĽM��@��ǐy��-I2㰳fy��&��u��1
�N���5�^�2y�D'`���6���|�Z��6J�K�ͻ��l�W�Hq�~|�Q�6[�E
��8A����S"Y��H�l�(H�	���,�d"�D�+��Δ?3P�0��@�&%�PA��P���&/,8����/�"�_t=��9���nl%Aȳ�-\hl�ɁP,���S��k�kU��ϣDZAk-�"�yT�����Ϲ	A��
w����a�ψY�śJNz��>�a(i���[��6X�g�q XlxVHYEB    5cad     f00�I3�9�]��<zx�1�(�#�0��sa*�l8`�炝��o��� ���"����j��p@���.��^�N�ѽP����/@ui�Ö�M�M����֫��J͙�tLW`FK9y���\ܴY��G!�<α �	�F�~��Z��{���0gT͞]�X����=ɰɀ�D6�ҩ���q_UםU�z4hQ[n����9�̘j]�q4�G�"���ٓD#��qHD�5�����X.�,��^ $!0����t��U7R��� ���ކ�9�;(�\���6��un���������k�k����iJ��Pll�=w\B��*�Qg�i��'.}���:�%�����kL'N�����R�h�՞�UDk%�|�1����I�p8w|$��C�7�pN�5dWĸ��[<{6d�����,�XR����X��\4=ޟ����f������f*K+�p%%f���9O�G[M �(:Ĺ�z��!��M.�s��4�mM�q����m�g:$���Adi��,/&��ZiGMiPH�{�z�>i�ʯ��{U�g��t e�R_�.�#p���0�Db+�.K2.7����rY��S�Z�c2�^���m�)����O�T�2�z���ڐ~����n$�#Bv�w��<�g9�iI�����M�@���@_f�2�Ha~�W�֖������4'�����0t�1�zd=:V�j���큧ʆ$������,L;0;S_���u�����ʲ����x}^&�L.���saz|Y�I֠�r��7
�N���V�Q�%ؾ�UP�EC���!čC0+����#lFgC�����]����3�B���D�F�@gyp��=g]w>�!u��F�٬pQ��/T�p@�y@&��m,��V�0:�[6 ����3yP�疪'ӯG�- 
��'��Y��$a�ޕ k��"�}��L� �{3a%-����`�[_�[���g��^�l����Wbt��ʜ��h�B[S8����@Tջ��Ǐ��?)�-)�@
:C�G�NB�����2DJ)ĩ5?$tA��j�q�ja5��!�c���I�Y���9�����OU�ݏ.I��+�g�̄�`�<�)�a$�f7d��N���悾�'����d?G��N�>1�n���!�a3kZ��7kVIV��m)&>˞Z��/|�Z%������%�S��n�G�5d�~w�po҉�<$O4	�׀�䡈���P���(=�#g ��ڌ�rZ���3nl&x|�QA�G1&��� v�l�Mz�љ�q>�Q�Ƴ��L��ڜ��.%Z	|�&�wod4Cm�F��H����p�c�����.C�E��j��H���'�A�i�]q��Z�Y囊���r<ݩ��%�Gy����ޖ_P�z���"�h��\w�]
ԍ�h�%��m���|+���X�"
�-:��'z[��H�f$�i�PV����X>�V���yr��Vb�'>-M���]9������CΊ�����jo�oCF���f�y�
_I��t����ڣ�ل��̈́��v9�,�	f1a���T����WM�B����D�<��N�DN�؀v3ӿ7*���7�>Ŕ�W��!�vCRTE�ǎ��[��/,8Pu�{b�� E}�t�W&�T��!`m(#UZc��FS��F,4���b��ݧ���O8�4ۗ
����S�Y�_��}vklӬ���݆��d}aW?�ޘX�a��;��14"�x�(�)��k[s��}X�R�i>�"a�F�1ù�Q)>FǇ$��ؙ;���ͬ�-�ap�~酄��xD��9�ts�^K�f{%�}���6����䃝X�5a*�H�
j��>t�1��_� m���{�޿
A��đ�C���F��w%S`7���L�?v�_o_��3����d3'}g'��ɀ
X*d�K�/�=�������<u�@ǻC<2�W���#xy
s�k')ؖv�2�r�G��Z�B
4zQn:�№�?�i�c��E I2�+�0E�T�2g�l�t�x��k�̗}ww"D����i�|~��b�~So��K����ѱ�.��}n���u��*��{N�/uA�|u�a���H2��KR8~��^F����F�/y�hNwm;�Q�S�dт��)���%/����_���bʹG�$�>����������,Q�W��:�؛�(gxYO��#)v�3PS���E�StLV�Nǫ��f�ݐ�������-��rJ%��t�7;+L^P�G�f"m`4�'�L�m��R�!�a��f�H64 �$�[�F@�H	��x�_G�j�J<���s������eI]�v8��Q�~�rM�~Ev�-��60@�5�׍D<�vPpN}ZI�nR����n�P�)�ͻ�����B�[>>�j��KFQ��[��o|������lU ���a� ���RK#�YAn�$��%
��r�j:@G�DD��g�f�}t\���!�{��� })s�_�M�_�� .e�!�L��f�q3�"[�7�Z�����yZ��f���/k�tMo���
{�,k��π~1ga%��r,Y�̩�˶�gF�˔t����E���$�O�_���8�.@ ;cC����BZ_���j�1M�������^�{*�S9^8G����y&�	d|u��\4.|)�A�Í�5p�����������q��,r wn���h�G�%���v��p���}����O���3mA�;3�+�r���9C4� d�o�i���k=�\�BA�mF��J����Cl����c�[EyB{�i���U���J	(7�LK_��x�����]dP�s`��G�h�k�P�O'*!˻�U�@U��.�֖v(P���@�\ؽ̏d�KO �p=����.���f���Ԥ��%����6����7a��/�9ҕ��{���A�d�UVWG�#P3�Z���L�QB�hz���W�����|�M\��^sc�A���ۊ!�a�i�A�m-k�����A'�	T9�:hF��\�O>0�I�E�Ȱ�c��ݵL�P~V�O�y��,ב���к�[�ֶ��_����K��Z�2c��Lmx:����ƛ�ݐU�_�*�f?4��\ ���e{e�{�eދ��o�rN'u��eǉH���2n�Ǝ{��w�@�~��w
y�E��X�+����1���[W����D����ܘ� Ur��>e�m�*Ze�^W�AI��u�D/�I�:��N�j�R��x��T>2F$5[Bܚ`%�����A/�B�\n*��(�I4�Z��u0&�L��A��yWzS�	�Ef�t0,fr��~���\��� f�8���� hK�b$Isd�X'�'���(�0��Z\0t7����?��H��'W5-@���eW�8���AyI��@���fIT>:z���7ބ{C&�fK`�ބG2�� �v�9P,�l\�bк#��� 53�O����� #F93̢���.ku��[��^���t��(���C�����N��<��Z��ې���k���N�"Q�����-P7�5U�/Eo�WOa�W��W�&�� w��zy�X�oH��"&���ԣ]���ZxU��ʖ �z�(v�(�^��k�%R�u#��b@dZ���NG"�S��J
'�T�g��׃�DA<P�ˢ��T
�S��h*J�5�u�����W�|��O��_7�E9]�ؒ��2�J�I���؂.�}�wZ��Z&yn���$)�jN��A}����"`o?ߘ������d�E��� }L\��"D1�>�W�y9�8��r0�=xCA�