XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ݕěy��+���]����J&?�eƲ���D���kY�p+ȱ�x*�I��FH��k�2B*� �fX��n>n�/��TM,�^^u�SS�����]��.����Da�v �'�ŢY�T��e���ٹ����J ��qa#�ԃ$j���[��ΩKX�k���� u���[(�W������4��KW��� �	ա��(F��&5�Ȋ����ֶt�\��b�6��v���_f����k�Ϧ��6W�(���gP��vN^}������7�'e�e)��$�"�y�)�o(}�Y��C;�[�\���\��g�v-�Dgin`{��ݙ���Ԧ){��ʕ>�]0ťޑ�Qb��j�3K�'�%����g��ێ�cAO���#Ɏ9٩]{Z������_����YQ�d���;!A�Dq�{��:uluX��Y�� J�D{|N7y�W]� %8}��Q��a��`�T޻�M ڻ<�_��>S���*汐+;H�SԊ!�f;��N`�	�[�&�
m������>���_Dn޿��"U�h�y]&�f>0v^^���R���d&��o� AQ��Ɩ�%��@�:��98�dѥq�	��DE���dl���pn,r��Dk/�*k8�V��5��r�܇M����'>�d��i���5G�!�9�̹�J�"��|C#I�	��]��MB��y�:������{�J|���qo�7Ү,�]g��W;73B�z�װZ�p5�x��1�XlxVHYEB    6315    1790woK�~�ў2H�o?�$�%��9�6�N������8᣸;��S�M��^jŠ9#KZ,�vpϜ/2�t.q�V<�n<�jȡ�~�'��6b�`C��4���W�)R?�G��B���f��T#Ύ�N��_�rIb�~�
un��6S��R£1���t_������CY���$����H�J�E�*��>qrx���A�Ug"��ccN�����j�� iֱ˒��N���LQ3��o���N����s�*멊qu�I�C��iH��3R�hS!��~1��x2��ĸ(u�3���p��#>�������,a���oƖ�-��ހx����e�Ůkҵx�\��$#~��!0C|F���"�Ȕ��/����bgQ��<8Ke�rykL�DHT�|�h.C"�%�IF[*��KW+H�쇹wE��F����U'o"�cXk�x(��?�K;3��=��S�u ��M�h4�0�t��-��R���T���U
@W�fu⪎�+_ab�A���{�v��tJ���5��������k�
�ĠFZ���t�sG`��@�G���5wg��X����W����P���jT����E�J_�4v�l��!r�?[�%��5��I�|�j��5��ȼc�Ӿ)p��;�!4��֚��9���K� ��7�A�Y�)��	0a�<L�@Z:A� ��Vf۝Q>+�t�k5m0¦���)\�l��R� ��:��9�Yz'#�!��B��0�3H��U,:������c%Q�q:o��ېa�v������_�Xz"P.�W���&�;��8	�c�_�.�Aհ��|�~�j�&D.���%+'uY�g4�űN��j#����1�ߴ�}z� �����av5�kK��G���F6� Duʨ�j9�\�=�sM��C�OL�?.�Qx>C��#����l����77���lf:��)�I���t�wadgD܈2�eL�;�۬���1�ig@8щ`ja���<i��� �����m+��A��F5�fȴ2\:�C�[����� &8�!9�":����ԗB�'d��AE�.���t�1��>i����繓�ژ{��9:��;���$="B��fx�50E�x-8w)�! 򈁢�:"�'��'�5��_�+�'�+cM��BB�l��b�n�9�мr��������"wA�a��@�I�%�sNR�1��!_Lh�m�]�S��i���p8r����r�l� f��k�M��������]����2����U�@g�ʵ/YH�q̜ŕ�A� �e	��4��JY֕#U�X`��(����rdt����j�lz���;а<:i{��L��崓�g�����@v��u�=R��>���r����0n�#�db���.g�#yկ7�8�}>|P��_�����+`�Ŀ>s
}!���p� چ|"��)Wݝ[�6���ܿ��c���C{nO�D|G�i��
���S��ߤ�Nϔ^
6��v�Zð��r6.4���=�˥�n�]�5�4�s��
+0{6��j�V���O��<Iɿ�,b����!ÙLۆ�z�?7ByNџ�j��ctu��~ ���%���S�;U�`�z�k�^Xr�iA,rW�1}����Fc����)�lBK�nHFR��0�+���uf�"�A��-�������#����5��L7��L\FL�Y8.�xn�W�m18���f�o�&�F}�9*f�e6�'� �sTN�_�-g����-��iFZ��;u�Uͱ�SZ	u�c���(��|�
lk|��=�p����o�)":pq;��QZ7�Î�A�q���!��D78���UЩ�n�$�팯���RP�p��M�\���'�q^�5\�r��v���'��:�	Y�O2��g�������߁�ݕ����׶>�8�D���۲z�`�9��`��D<)U"��Ssx����1�н� �	��I�-�k\-�V��Db���V�[ �"��@��A�{�|q�S&�RnT�� u\� ��U�L!��K�՟���]�Fe�y�x���2[t�|e��mԲ��G8CC6�w�'
-o���S�o8<{�cY�0|E�R��&::��Z�:K����v���1.���:e�ӭ	J��v�N�2��C�y�n�-{��>�mk.bg9� !���U�}ߡT�]G��[v���Ls��-���)�I^ݪ�G�Y~gx�@����S��6���\'�;�	�x�v���~�þ�f�07LN	f/�{M�SЈ����|��[ҍT=��}�l 9Lx���e�=X�9ؓ-%�!�~_zC;����Vih��M-(X�Cs����DDn�*$�^(�Ǔ�7���|���yD˨��9�K��w�NI�b��V�Ɛ��о���2�ِWG�`�8}�p�jgGO?%�����]��i�mV�Iv�R/R+�N��Hd֞�D?n/�m���[�x�U�3֙��*H�̅���<�v��� },����]�T�X��U�������y ����lY�%н�[���W�L��2�"�Tc���i����������ll��P}�2|��"��u�8(����U	�����_bM,%�SYx��j�����LV���<٪��]�*�@r>� ~z�p���𽕒.�D5��n
8���S�6��JRa8���.6���C��'�N���o�=��?�%��m{�K���a�k��~;:��e�����K+t�>�1mZ	d`L*n͑b=-����i\R�S�9�w:G�iG���٢��� �
�y�g�7���/���o�%28�븧��d�!�����g5\��;p�xeD�y��/���G��o��,^F���1o�XG�?���RE>��TuNڼ��S6D��*ؗҼ(E����
���B�o�"i�ۀ�� ��b����t�o���9l.��V3PA�R'��32��H����8�s۾
߾���Ö�70�|N��j�L&�_�#$�.�.��[�2Ʒ����i��5�#�y��d�$�v��wD�`n�r��!��H��<���S-ί�#�cOC���\d�=R�¡~�F2��Fk����3�W��[������7����![�@��Y˥ݎ���2�w�}T�ɕ�ɠvH=g#�P�0� hJ��xC�tT��E2-����3�	�AMi��&�Ӟ�BZ�D�<��s��z�_�! ���F|�x����-�`�ޖpP|fZ��"2����	���涠��Y���v�
�"����PMEV���	����2���N�^k�/�������%G�V;�?�J(H*i���bH����ȴ�CB�Jn;��o_Rs"������+�Ac<��H����Ӥ`�|1�8��3#)��<���S�k�ی�'�������&���*�8s�h��M�Bh��QO	�Pc���W+p۶$+�(��R32���&��t���� �]dQ{�^��+���X�)��f�З�md��)欭vƍ�\Ν
n8������߫��?� ����A�s���f�m��&��F�ɩ������̶����e�J�_�,ZAzj_� �s�ǳ��Fȑ�UNp����Ú�d��Շ�ò�k��y��M���J�
'��3�P��#ʁ.��/giw�FJII���Px�SO�>�9: L=���������[Rc�`�R��@v��RJ�Re�Ve}���䚘� ��=���ED/�z"%��9�RYz��Fb� �Է�t�;+6v�)�}+��Gv��}nt�k���Y���_��c�������ݖX�������B. �߼�l���8X7({Ţ���6~ƙ�@rδ-���_�������\-ʆ����]>d���g<�a?�J��,xd�Ӌ�d��	F�u���u���\�1l�s�Q��r��znC��}:��,��ijwaϒ)@����8T�%�>��ݳ�����^x ��×�-�@���%+ta�ֲ~;"#V���4.]ΠExuM�?VL�/֝����)��r�ofD_���7�F5� a�6�C��{8��D�Uu?߇X���՘��)�Ns��[�'�zڕ��PH�`��۠��F�X[�Y�-�2g?0�D3��&��J�j���V!hgg��Ϳ͍�T�h�.�3W�:�$J�E�JG��/�ҟx�Z6j�u����7�-%�
h.Bo�}�A1{nH��@�{�y��ݣ�tn�)��Gn���y��3"�D��T�!�h_n��!����_��q���7'���͋U=8�ߣ�fө8+�(
����q���Uu؄�̲�g����x ad;�~ˎ�=��KX���`�;Tq'�ma��\��o]���5+K�bu\���K��-ʸ�eUw�$2�ڿ�~P� ���į�\�X����<�N���i��c27%֢(�����^�5>p3���)��	�#�(`��1ȵ�佽�B��kS˲�4P:��g6F-m�s����^H*r�����Bb�V�t�~��w��Rw�iC/�G��6�
Ta�HE�Bgv�R�9�����V_=In/j�7���e���>AC@m]ΑS���.����V�^�ifw>�?k �z�NGs�t�s�mE�?�$+
^V���[�0r���G��e��h� �#�h��[h�i��Fu��;RY�ʘ�Z(:0W��r��qQd�&�˥���zL��y|���/mN-�&��2�t�1Tޛ��sH�i+!� ��L�=�s��&�kmb����~�>L��@���k0(y�.�i��p�%Nҥ��w���NL6�	��_N� ��x<k��2��4tg�G_V�՚��V���$�;��x��`,�ǳ�1.w���8�=ҰX*	���+�i3[՟�k��Z�"97|JCy���Ať��d��y4�ށO�1�f�:�+8�,��� 1���@�����Ys���D���H�߇)k}��ֹ���Pe���=��{ܷ��1�w��F>�D%�ڌ��mI���>hS�^S�h�i#�qz�>/� �Ρ�Rp����$���%�{np����ΟRQ/a�3]�*��9Nc� z:��Eԛ�vE��y�ORvN3�7��{�-�3��K0�:�%d�}"ϻ�������4ԡ풍 t{�m"azuЛ�s�(�!�9[��x�z�xw9�U�V���ǀ���~���,�Q�qQ�o�c���uP{\K�S�,A�X{�0s|��"u��=sh�o5
gXNR?$�w��5�t�M���f<��D�5��<�]�	Ӎ�L����"�MJp��[�L>�zED{Y	Qc��s�i�hV=��[��=N��Jb)�!��.Uf�������H(��K�C۸���_��9c/��s�D1%V\�,;�1~}��^yh�%B.�,em�;QK#�*7�7�릦�'U�G�wr�f��!Tގ�a]��Jcͳ�Г�Go�����	n4LnZ�h������?�6���H�t�9|Jv9[�T��wb�,�e�����_^��)���*E�����o3t�&��v��d��^)���W8$QٻK���D���F3����L(����a߀`c��2Y�Mxa�2�.e�P��}�%�;������NH���~]r�_��U��L�HA��/a�fԪ�b��.>�� �R�.���]��C��H�n�4n�d}��?c׿2��N3fu"U�������a���~��&t�v��_�k�[�sc0�����_r?5n���%mT��p=�X4�BV7kWy�VG�D��Y>!Y�-�$6�C�Y�����ZZ~˔,6Q�t��zd�̫����M��&�@-=ƃn�1�YWp�`<f��#����q86/�����T�[C��7AVJ���䓎�z�;�_�f��������1��Ko�>��_@Q�H;�A�}�]I�#j�����~w-�������眝