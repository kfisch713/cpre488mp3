XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��<53�Χ�c� z�/��%eN�q`
�w���P�m�aF� k���NE�a&YC��z�W� ���[x��0�u]�Jh4pS�N}w��0�m����/��kR�V�Ac`�������K�ǑY��s����3�R����v�Pa��nR^�����{�XR��&�DH�eêt�ep�X��r��+哟��,
��/!��i'�cϻ'$	�T?M 6��%�`����oK�wɳ��E9b�i�oSopgm�&�"��@���!lz	�ɺ$����b'���0�~3ܦ�WD�ʴ+������z��w�;�G$�E@Su<�}�Z	/~]�LbU���-
%��:c��B���M���R�>R�ZC����CG���W
�ޡ�Q7�����Ï�-�"[B5��۵S�uص�}�7���P�6����`�_O�
��b&�N-n XZP�|����N	�q_>φ�k�|j���i#��-P0;������?�XF��z�}�)�AZ�ǩO���~!@S�6S�����W���pע��V�3�8*�6x��!��~-����,��[�I��飔���87�N�T��|��.ո�\?q�x�@cH$�ҝ�b���
Yw-��S����i�&39ɻh@ͣF
A��D� hU^Ѯ^��7vH�$g���S��e�v����bك'oU�1��v�Yj^i,���Q��l��U&FQK0`�_x�������rY�Ц�7
���F���	��x��G��>��f��řXlxVHYEB    fa00    26e0)�o`�Uo�MU��J�)A���&^`,�=!�E�-Y���i;"����2D���5ߧ�`[�� ����R�{��vp}�0Ve���#����F���Dz)�z��J��m(g����g�&r�|����vg�^��O�˽�\Ĉ�N��k��{�0a�KGL������7���O}�u<� ���*���?50mtR	�4�sC/"�8���V���_	�t�0�ՒWF#���9�W5������~�������ʂ$>��e!R!��72���B���]t����� Y���j�����G�T�4�^Uυ$��d�h�{��7և���_0�̯�nG��3(W>{B<㿈���-*���}3�c���OƦ8~X��Ƨ*��nY�U�+R,�-,a���s�����Kzl��&U43'Dq�Ñ��ړ�>�i1�[���r�)�k��C]*�����]�xG��l�g��V���ǈ��|��;V�f���C~C�G�ܐiW��*\ ��\M[�h�A:OLǸ2"0���U��OFS�ki�M1��Z����8�{���2v?g�:va�*
��5Tq��17����nf�It~o� :�o��g9�I��'�\W�Yv����w����^�R�k��i�-=�\�;����]�%p9Hu��n��	�U�]-����bN]"������wb�f���u���d��عg*�������ɭ	���)�W pG!u��,�V��^}7챐��qT�r���2O�{9���0�pj��[���a�H�'�SP�9����ӓ�BR��I?�_%�宜��6P���>���3����HF�w��0�,�Ƭ�X�RWyP��\��7e?֎��H�綪"�>�Z��`� `r��.̮�|O��v��%Q }���'�0���b��I�I�8�Q
N���]�u®(L��aX+�v)���n϶��T�b��q�?Ȣ���7G��rr܉�0ڥ��T�A&F��,�5�x� 3�&�Y_1�z}�"ɥ�Y�N^�?{�J���'�H�I5#�
�ꖶ^d�j)K�;���j7� ��GM�N�f��Bt�q��G�5PҬR��V��N3pU6��f	�L���O6��
K$�4����!�
��7F��ǻ!���~U�\�����Ց��gƪ��\�Ł���_�W��Y���Px�8��M��~P�\���h�g��ج���L��~۝��W��-�3�v�P'���a���Y$ϘkIk���k�q���,�܉UA���t��ݨ@�B�Z<!��c"�L��;=�ѐv7(����-լ�K�'q��'���L�z��}���%�����|	k(�$@HwK��Bjm������I�5:xe^���~�ౝ:ŝ�!�8�#�dc:_�i��s��y �ks�[��RƸag�%$D�Y͠��_y�㈖�)*;,D�/���T %d��޴U!���농Ӑ��uU��WK9�_�Y��)ҕA��x�TR�׎�J��,ѽ�z̦�i%.y��@6�_�{��D�)�'�	ڎ�E%�7zv�R���n~�"=�i�0fX�;�8�8 7�xP�1k.���>�i\�1*x9;��������%ĝ=9P��L��,c����ݏ�}�&�u��7����]~v�h��o&�X�v��^oI/��7�#�D ��ι�I
�_v�������s�u�8�lm8<����g��FY�x4����/y�sn�^���Fa?�G�~B��:�Ww�s�܏�+��]�lkI����~�Ea��1�����H�)JZ|��cZ��A��cR$�q�Ƃn���W}"\�f��%,�	j�뻨��H���\#
���4�V���w{��p��h�5n���PD��y'N�A�;�Do��w� h2F���HգA��зǓz�;N�Q�q3��HՆ���qZSʤ1��|��_:s��X�r�R:��MUԈd}�׌V�ā����+!\�zf���v�A�q4�q &�Zm�[�Y��*VKj'e��s�/| ������EꙤ2�}��8M�w�W�<�)	e���*v#���Lc����W��(ɱ��ׁ]�eA/��a>(U�-Qe�+$�� �c!3�6�j�=:����)9�q� s���x-\�D�V�[ַ4U�K3e`E���\ [E���%︉��M@��)���~E֘��H��1@��*g5M_6�P�*��Ʉkq����4j�`)B�Hs5Bs��xK;-{��`{BFo(_Z��B�t���Ck�x��`���WGY}�H�>:�rD:49ㄉ(�<A��r�)����7�x���7���M4�BU;U`�D��,饊ޣVa��Ň�[S���<BG�{����̠�	4����jF9#��HG�v�EUhg.���F/�%JƲz��5�0}�֕	���	u������?�8�G��P�m���Ĺ=yk�6n��͗�^������i��!nu�M�a>^�£?n;g�zz�u��Y��� �(�&M����j�/V�@�Y���f�i#����l�>B��4�������&c�Ԧվ
'�
rxg�K��_�bf��Arɵ���/��[�3\��a�'�6����,}s�#رO�����Q޵Ò���4 !��
�#��/ ������t�� �*X�̷6��iҫQ,���so�[��ǝ����8�r�����kAjH�`9{?�'���ԶS%s��]�����7��*�f?�[��yOhm>9�Ӗ��+/��r;�Tf�[�4"]��R6�B��E�h)!��c/�D���$\$b�'�m��\n�r16��_��iy��E�I= ���p����P�&#m������~�kd��?�?~Y��R+��Y��0��ES:���D���!o !��~8��o��+��1�OƤ�N�`ZF�}�����[�#� g�Fi=/	�ʹ�V��Tî��ъ�o��P"�h��&�='��c�r��j��Y�2sј�\�#�k���I��e.�Z{$NߛVkp�߿��Bx�,L$��7`75ֲuے�����1q�jk@Nv�!1 �&3�m�.��&CV��Wf$Q�[f���$G���B�7�U\�<�^�8�X�MzM�b�8p^�[�����:�E,��+�wm�%%tré9����{�����>蛿�x`tѭ����zE��~�����yq�1b��,���FXJ�ޘ�&��p�˫Ѭvh88��X�Z�[9zއ��sf�K�^�R�� 2�j��bf��V�&�9<3�3�-ag��`~����YA>���E�~�[rU�ۘ�GN��9���"�dxP��Wk���T���.\ h�ҿ�}#�Z��`ݺ��3�1��)(���q�	�_�������R���V/�>��x9:O��HK�`ɩf-*����R�/��5_ۺAg�Y�1R��Q�H��ھt�z˲�v=���N�Dps�V�%�|eC"�Ou��7xU��R�>u[���+�V����<<��u}I�ӿww������6���� ���[ζ������ӣ[��})B�NW��
�P@ ��'�&"�Xy-��/�B�K���,ヺ��zk�s��o��]��&W��8�d*�FhD�*`})7��=�~~y�@'F��j:"�,d5y	En�%���q�=��F�<����A���ً׸�s�D����{�1��sM���xO�2�˨��i������r�^Yx{�sT�=�6��.`JU/��$�	jhZ��Y��D���E�aBO�;T0�q��s��l��=�o&L���3�8-�@�)(�Z�4ڎ��U���
?!�.�Ӫ����q�ɿp�tf$�O��.�*q�RaکH&��~��4�1Um��?ӛD'��`���G�/�[�%>�om�\�oGl	=���G�=�X�R��*���ݼ�8�%���� F�+�.}�	���ΰ� 7� �����U8���a����o7H��j4[X	�Hf�*7T!@4����q�IoeH&ٌ��fa��ݬ xo:� [�F��9��|��E��y���L�wI uư�μ`Tᔍ�IV)�U!�/R�%�
@~3x;��+�ڎ�Y}yy���3(id�zr3��~9��)���K�0�ͻ9�b�ڠ�V.r�v�#u��Zg�q�{��W�8+��gA�S�b����v_e���Q�ս�W"�H(�����UK��#�ך����;ڛ�U��E4#:���� D���	�[8�����Ǯ�\md���U��|j�@7̻�w8-phm��ʡ�|KĴ؉�:�!rݨ�����F{�f�Z��+�6���Z�O�j�P����BB�@	/UB�f���x}��Ìh.܈��YX���n�\� �&����G;���$��i��� ���cB���Ȣ=e�������e1�;^`���d����=��3��}a�����!��ƹ�(I�ǀ#�*�x�����%6��A�ނ�-�6�g��AB�_��W��  |_��F�x%l"�8q�
1����L6�١���#�WL���]����VP):c�~���6�J}�,��f�؝o�h�����'K���%/[�X���}�`a;����Jo���pa2/��z�2�g���iѰj���;U
���`��|؋�
q���wyծ(5����y$8�p!a
)���v�v��P {	!u���0�Pнw��P�(F|߲~�����|��wp�;�$�Ӆ��ޙćkiB�%<N�P[����F����<��CN�D!r��Ȱ^c�Ǹ&� �DΠ�����zsz�#`n�л.�ʲB����ɨ���mZj�nD�!��l>|��`�"���E��C$>�tL�=!�ui|?9t�)�+r@Bnt�D5>-cY�����ڕ60� Y��=:�AŴ"N\�q�(�� ��C�ex��T�=8:�PDᦍ\����g�.ǲ�����^PU��y������RZH0"��ߠ��t� ��S��RH󡘹5�A��"�^.[L�	���h�7��+��R��S}=�Qŀ�2g��ϓiBQ�qu;���R(�ŖSSVK�|F��ic���	�q�,������ǵ&q�P�#4��z���Q���̪C>��{U:A'���
J�~�ٲ�?���
@����Z`����j ������ $lצ; d���'�,4�7��b6��0��P|c�Z����Vy�Sd�Z�u��6�A׎Z�-g���@�ʋ�4��X�(��n��C�Ӏ����鎢u�c*�UwJ_��hKc��v�����Z�^��ߞ�M'65�\���F	�i,Bΐs^����Sp�6�o���a��T�juM�GP�@���`N����8�i.L�kԊȖI5:_qg֜������A�Q���<=�V[�7�BGx<���h���R(uA�:B8�/�y�s k� ܓ_[_��x���6գ�)���Y�]��p�6���S#f�Za]�K�cd���h��K$�l\���'p:�o�|�o��y�����2KA��:Gh\ �#jk�h�d��3%�̴$��O���=�^�h��*������8�Jcߏ�W:���:����ӵ���/\��v���k�nCǦw���9��aV��M�50�0�4����d�dm��%w�}@�s�Zwn�8�%���D���M�2�����q�1#��NJ�#zJ��<8j�h;�|�X�1�Yß́=+~���j���̏���X�!{�?�D��f��o���zaE��:-?^���O�d�U�r�/\�Jd�ۙ��� 1f3�5�p O����:�̨��{�
���������hT���ѱ�C����!�)^���~�v� �hP�w�[]:/At2Z�eݐ����!,4�Hʋ�9���d�w�0�����.��N� ��%��y�<�K��|�R���9���%ka����n:߫��h1��c�d&�.��o�|3;�L�c�c�{����^�H�-�.VB����`T3+^n�=��"3C�x����pf}� �,�od�SR0�ƪ�:��U����ݐ�i��ҋ@�����}%�$2#���{QE�J5�S�q�:����[��>p%�d׈�lP��4���`ΘYsT6��B�ra�н����+.�qYo˸��2�y��w����U*��מ�킆���&�B�F�`vV0�iyc�lHX����ٽ��'�R�h�Os@�&��c�B5ԉ!29 �~DX�s+%�-�O/UT>Ό��T���.�|6QA*�6E�1��㣗Nru��pR#iv��ƭ��g�"Mf��H�B��5#��˫b�y���|)z����
<�Vm%?XiQ�A�<ϺV+�_h
��i.5��
��� $sj��T��ǣS�]��V��*�˚�}�/6/�=��lV3k��"��:��Ӊ�!73�=*j$S{[�Ul�μ��)��� �of�>T������ލ�Rv�`Q�s7��Ҏ�?�����7N~/W�����
y_��]c�A�bG��g���[P �`ZI׀���_���Ǜ����kA����~��VFEX-%�`ͪ�(����A�A����Y�"���{6��S�*���܄���|ҪN���)0F���V��m�$
l���Q2s���Ђ��Pu���p����&������'�\�cJM6��l4�N"ߗʵ�;̚�)�`Q�C�f��z�:mN�?H����-����������,�yc��Y�z�*`��}`��I�VU�����5oe��E��t�e��_�q�G��M�2�&]�������B���a{_�h��?5u4�q�|Ɔ~��$.:��:z�i 4�5o�[����H����çxE'ƹ���HlA�b�L��W�lnaY���}Gè�ix�ˏ�= �����!�0�ab�yC�����!l��1F�Y�[����cX3 ��G_�:9���P徑ۏ0qdyƃ��?n�F��s}�&������&��>�/?o�� %�U-XޙF(@i%�����<iz�n��)�8�7�^�H>�0�dy���t�$����W"�Դp��@�h�?WX����TH0�@+��<q}�oȞh�ykz�1��T��k�ErI�p��u#)!�F�X$�!��a<�1��ׇ����X���,]DV�c�L��3ǟ�(�1��))z���Ö�i�ʤR�TY�P��taZ�yk�w�����)�`�¦$jY��.������g�=J�b��L=yM�F�ڮ+�ԭ��L��֙.ΡErElC#���/'�޵�@�&����\M%�CN�f����n��/yEU
�$��$�E=�[.b���7�>�H���8ǉe�|��tD��~G��y���ddN�y�ڌ�7���W�h~����7]���o��>�f�c�8�Kd��6�d�x�s6ũ���'�D��E�$�T+�f�ǷV7�9h���v��g�B/xk�y^�	+�p-f��i�/��lW�	�S���bBt&�T�A�!iĽ�-�&��:�!1h��ˀ���;kh�c��p��������=�����I�I��_x�_�z�<���=j����r�9�th�D�kO�m��_|a��BZ8�=����I/���~[�]�ݛg�=��e�Uu� �ur����6јtX���ϓ���C��_�{�����g\Sȥ/��dr�4�n<|��U96�H��GR�$�X⾞��Ǳ�M�
����ت#H����%A�3����l�;<ߨ���{qI��/��ې�i�ex�K�pg��_j�F<��r;�r�#|
��°���=w<^kd�s.ȻW��>��*GM)7��j�?v��0U#[�xB�<uO��g[ΊP�ړ��i�3���)�B�\�;�}3���V�?|�{�>X[��ǽ�V`$)|�y�i��-n\���sȔ�"�`�fE4i��2��f1��Y��e�tpHf$E�|㱯���(����p�A���:�uuY���؛^Gۍ�a��ײ�y]n�T�#�9:F��Ƙ��_����!x9"s}�cN f��!�:��e�f%.��ELG��p}�5��Ф7� ��
���9�� �&)
�$�K�����q_���D!���P����fl���p[V�L����I&�ك��S�z�B����Fw_��P6
Y0�u�UakX���'��rJ�֦/���9�P�������-m%�m�K� �����ޘ���-�e D��L��� �֍�g�c��rdI��n{r�X��t�n����������������&�T�Q
��	����9�K,���1�ݨ!C#� A�If!�EE'�c��@u}�����]'�b��
�(�\�4����%��7��BZ���S���X�t�a�Z��� ��pyT��.���[�8.�Eq�k-s�.cܠ�v�Х*��e������ ���*�4�z܍����l%��4�gs�{���YY���0����-�.��U|�[��
�6�"�!��5ه.�\�k��@���x�!�ϕ����7��W�>�����~��AJ8#���{
ݔ� LФ��?x���^=���qT���h(�)��-���Ԣ`�d�n��t�8q��`0;�'ɧ�w����D9ν��s�c',h�u~Yd�i��j7�l��<��p'g�2#�X.��z��K��	/��Aִ��>2P�M��} l�~��`3}��}�����H��P#�����n�>��c�*c�if�.F��T��M��ӳI!dJL�K�`��s���{�^.�8z������\z�� Ġf@w�N�م�ȣr(�&��R-`RP���S���ͷ]�U�͙w� )7h��c3'�TF]����q�Cw��0C�Ux��9��r�1&�,_Ceu�@��q䣷|+���q��a�x�V�Gx����w�SD,��;�1���A�y2��,,���뙯���q)��L�$���(T$��ʷIB�C5d'pChW����z��xd�%q��ꊿ˲� ER�?�*�к��ɔ/-4:�m���C�?�Sқ�E��~��WI^ .8�M�]�% &Y��w��^�����g�׍~�͠��1Y�b ����px��=�f��c�|\P5��P�RGU���Uy��$����=_��V���̄�CMs�!�L���CwrK�̄�d�s`�X[��{�V�H�3߿`W];b�p��qG"5�a1��e8q��K�G�£8gW9<���.��c@���Ё\h��$��������S6J��+Z0c��m�Z��N�`��6��ax?WK��?�{�x߿���	쀈����Q\���m�D0�p�ݬ�Mǩd����Ѹ9�g��iX/;UW�I�Ȑ���W��8�� )@H�t��l�}$A8G��>��6�^��&��LV�,5�d�?�m�7D0LGy��D_�1t��N� ���'���S���)��!/�0�j
�����n鎜*��F�Bw���8�|�b�<�b��i� ���#�����l�� ��H0��d-޸X�[|; GX$c�)�R� i���kGp}�-���L[k�+Zٳ|�֐:H<MX�"���j�'���`G��Ǘ�~�Z�lkΛ�
�#ۢl"^n"�}�b� +�m08x�0i�TD6��*1Zi���q��m��K��K�P��l��d�����OL�$5%�e~�֛�*ٜ��R�d��|c�B��J'�/P @ʢ��Σ{�c?8�J��=��>�c�)�t��
+5����������]��%��9�>�C�1>����D>�c��Գ�1��-�Y���:���́2�+�k�s_I���H�`�XlxVHYEB    7d55    1450��~G�DɐOk�,G�RJ�ߏ�$���nK��+��6�r��D�jo��g	��㳥�P����G�V%���'��vL��)򼫅h�8?�7b�7�n�C1�L�}��	}FЋ�Jz�	�+���u���3���m�����#1_���c��p�	Q]=�}A$X�V+%��/�y��7����Z�1h�/��[���gC��kߋb>8�p�������׺�A�DhU8�H�^W��9�W�!sgMq4%#4"�	&����"�^?�Q�8Tz��p>|�
��LJNwJu�C+A�_���/�#�8�ڃ�*hB��d�ֽ�][v8�Ol!'��7�S�QXH�hmj��s<PX$/��۝�k�x�O�[�SD�ʒcϣ��6����2����m�`���ͅK1	٠�=bT���z���:S��,��wv�oV-\GB|Îa2	aE!����=���+)������rx2'*fb?��K�׶[��O	���@���],q?x�b �͘'R�D�5���*k�?p6�k��i�	�ԡ%Z|�p������[���tBWe�R�T�d'�ƉE��2(2vK$�M?�7kAy��[�C�h�;>��p;�G� ��ם�Ƽ��6�k�=�uݹJ�PS< R��rf�`�v��,��*��y�}V��Hx�H.vX�o�*��驔ƻ�b��i��B���搵�Z����W�_�*���_�=��w`�lnG�������ݬH�n3��)5F�`Ksl9c	_]p����Ӯ��N3�� W6�O��H�8��ś�V�l�-5dʃ5k,�.ȇ4�<��;��ϧ�:�Q�jk�h2�d����"3��j��qmR�� ��;����rC9��V�'(�5���a�3�7���\F�T&l}�v�tD&5�k��Ǽ�Q;�%�]���"|b���i�����֏)�W�lס:���=A�q��{�d���E�I z�(���p�-�*3�r�OAM�2��t��lSc�����I7�T 8T0p�7�0@| Ǣ�)��p�+I6�Np����?�ɠz�����_&��Fv�+*�8:Df4�C)�Y��z~c�@�F�"��F�L	��,5����`�.�d9aK�-�b
�c�G���j}Kt���?�n��0����		�@�_����1������7�,�v�í?P�<����!�4�y��$Wڱ���yi��q��(Y���2�=t�Bn��վ����:ݭ,�R;C��O�ӿ��? �����,'�Zl�r�_�N�����xOΆ����d�>���l�D�A9��7��/�tP��R���GS��/�"p�@��y�bQծy�r�_5�_����d����t}i|m�?<ڛ~� �u�1q�D�|8U�cg���|�-��� �̚�_��鍽^���s!����v>5k)�a&�a�/o��:f��$�SK�ER��P���̶7��ei�7s��׉�jx�7�����JVNm5c۞�L����u�]y�����s&CJ�YK{�]���UHy=���G��2zN��̪�j��)?��5먃�	&�V����`>���l�cO���r��ǅާC�;��#J�y͜��R�f����\�y�3��R~��c������ꌪ���%�Y����ό�E"o\a酏�V�Y�9��1�� p���lؓ[@~�
D>Or٤s_lͲ���'P�G(��m��[:mߺ�H�Pk}��o��h}�?��>4G䑳���Ν��w���̉	:��Pקi�W8��Zb��oZF��,ox|���G}�B��>C)�HYp �b���$�$�x��#��@Kde���[�V�['�ۡ!�ә�F �O�H4{f��K5Ӫ�fN����������L��B���Ĥ�l6�L�U1��w�'�%m�?М�6�3�Pcy�±r��զ{j�-��0<	^b�"�sf�j�\~���x�������N)h3y�n�K�A�ڂ��_xiڇL#K������%w~}E����P�Tw,>K.v�@���Y��s{��J�RO�w`��@�. �� �'S��F��v}��P�u��e���1�}�,F](��i�G�_���N��-��\c?�H �V�ġ��s�Q��P�S�S7��cv�u�Z���j�C���Щ��
 ��1��خ� 	�hc������M_B�Ӎ{#Y�%�l�(Ћ��ik�.y���x�d��lx�z�z���$��Gg�L(?���R�Ƚ��_���O� ZQ�f����w���	�]�Ii�r�p�c:擦/J�\���X��IMj�a4��Hb)��>�`f9���t�p�ҋ_��쮞�i��2:ѣ�
<�9��C�Q��s�������Pɺ�_���#����~��0kM	j�N$	� ��s����s[Z$�Y;��ڰ��^)!�K�-���Q8��g�^ϖa�Li��p���%��xU�����?�(���C���{�Ԗ��猽=� m$`�����������_�������C��ʛQ���1LbbΊ�&��ӽhUR�T��\UY���DE���6|�M,V�L��x��}&I�Q:��ėMD���O#�i­fFꂖXF��7���d�-Ck�Htd���D;��ߥ{�?���j��*P�ҭ��׈�!a@Oùe�}|�@�-��Ye*��?B��3�'_�-\3��O�������t#%�gN�=q-���Ty�Ʋ�+��B��Qk���_���w�[]ۣ+�h(	$�f�ҝ-�����=~���^��c��Α�'�d���e��7���o�W ���o���P�U�`�r�paTHS"|�[�FM�ip�xFM�p���R������^�H���}/GFH�>��c#?�����s�x�.��<�~��)�}]���%��(�@�nf�)p��`Y�<�U�j��Z���YO���Of��M;�9/@�B1^1��_�ǻ�߱n�6�ܾyZ��J�d�cӓ ]^Á:l﨤q*�:����	��ˈxt�ۆQI�V�5�����Z�Kh��f�����N�DR봅��~�;ǝӊcgbi����X.��2���w����${(nB���{����	vgm �������ɣ[Hzc	j���M��Ly���S�����JQS?;ˆ���N�H:�V]t��I_���^� *�U�%�ҝ�dԭ�R�?b���Xw�UX����0̬�P��Y��K���I��̇+n:�-E�X��� m컴�!����$+�m����0_Tg<t.�8�a����h-�3h
��!#eMF�]�v����Wg}�2/z�%;�x	��h��hl�~��P4Q�7v|7/*6�E�b̈́��T,���S<�",�+Q�6W6��x#�7�Y��P�C}Ydm9MҐ��F�O:qXW'���ڊS��~�l�I�Y�[R]h��-l1Te�6��g0�f�Q@jM�1�)\��a��c�~�(!+�:�_yH�N�>>>Y�����~c"����e{��8�?��緿b4���~��U�n��G#�=��1�F��b:�����ٌ�T�˅Qn�@�)Rj�
�x�ی��.w$������S��V �e��p%� M��ZI�R����k����D.����u�!K�5XAB�%��Z��
�x�Y���N�@*%4ʣ'AmF���誘��P���\&4�`1�D���S"v��)i��_8(�1�揯	>�����͝$�3��V�}������0>j�׾�0�5��5Z������/cU��jF;jO'���B��/�����òU�{�yU�,L�蟞��A~3߬��o`4f�X�5�T���t�"�e**�Gޜԧ]Y$���<��j�U�_��|�%+�U����IZ9��EP��R�#r�R^B}��8��"f��	�w@���vXҾ�J����������P?�ܷ�8I�)��hi�첾I�	���ۄ~���8�4!�'�|��E�~��E�f!�o��j!#�_�7�;b�,����\��8�N�ˬ*��o@|ܠ�fI��/%�d��VWWh��b��D�e�$v��

Y��e�Ϝ(���%)_S����$S����C'��P�?��{Kz���� �q�,Q}ׁ~��U�w�����b�c���"j8Us���r���-���3D�#��� �I��m�~�U F�a��Q@�K���vq��X�l���E~zӬ�9k�4� ���J�K���;z��e;�nQQ5ST��}�7��D3���Z��y�l��2CJ>��b�l��+���n��^��,X4b�Pd���WD �_dL����u�W�T�˼�`'�1�Y�)�� �Z�0O1Ԭu�T\�T�+U�N��ۇ�P��&lB.�c���?�5A�|�>�S'sxȡI��F<Ȣ�sҼs��7i�ϔn4K<��z���\s�"JZ�-0�O�֮}��g��{9�)L���KUTɱ�,�ۦq
b~��IW�(1�k�o�sG��G��|��pm@n�t2@���b�Ox^�\��m�ա�"ҋ� �G�5� W�Ӵ3Z�3P��;c���/�5��.D��:������m6�1MVۅ�p�ݰ.s506$�vr'8F�PW��L�^^�����k>^�%o&�e�TO��n��@�Y;4��i<�z$�C!�:�rL�/�EX��9�*߇�ުXk!�P���^)�;rc,�C�� ��� �L��M�m��W�����IK���o´g�m����.�'Q�{^��Ŗ�㞡��k$�s�W���\�;0��d PB�5~�NѶ3�������d�O#�s����Eo�]�Pn����$�3�R?�5#wK**�������)?�9��!lQ	�=5tN���ol��f"�0닚N�����c۸]����w���Y��C�n���\�uE��ut�ϧ�7I1�[ס��E�e(5�"w�Z"��6F�r�l�����!{���SO�����
�c6��а�1x�L$����ZtF(o���p5?!��%�6�ȹ̕:w# &Ʈr:��׍�f���˴l�� ��.��]��w�@�x6�JZ�dnz*�C0zz�Q�/і����P��@w