XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ڊ�O����v�i��Pbr˖��	�hY��˱�ۤ%��"���f�J��✋H�B��Dcԍ�<�����I;!"�)����(Y��<�I2�kF#a�x�3�i���_-"��~����.�ѭ$���4�ԖC��E���V��t�#
���P7v-��l����*�#���S�^�$j� �c�N ��jZ���1���ƔH����/Q~�5�J;�h�J
=SUչ���m��(�X��d��-�\H���M�d�{��+�d���j�Ȟ��Q/�n�oBܒͯ����l"�p��!������4�[@Y�<F��u]r-M�yt���<fhn�~շ���·�D�ĕ�����$�"v�Z��7��?�ϥhⲥ�����E�NJ��sO��z�F�;�M�G4��u�E����DG�O8��(D�e@��B<%q��?tx1�����c�8�o��-��#ò(�и�ԇ��آ���q.��^3k��W���VL۩�(a	����?�vќ�9�����k}�5��Ƚz-@V�	�Rl�yC1���{Q^Ȅ1�*w�x;�*�ӯ�a=~#b0M�pfS8ᑠ�L�'|eD[D�V��$�X�б�����h�!����g�Ή��)��ə���'�ⰅP9�j�#�k=l�:�1}�>�h5J�T��kG�i��;A���F�&D�cAd5�T���55�X�ȝ�m����t�%�@ť���DA>Q�nق��x���+�*�X�m1�Cl�������XlxVHYEB    1a34     990����{�7��%F%��z�h�;�?Ό���­�l������V�Eܥkα�~��.�b߲A�����EI��{�n&�n0���5���=��P kǮ3Z����\�$��n",$؇��¢uW$ݍ�D����ލ�\y��*E����u���������*����.�� F�����-�N�>�h})�����ٵ��Ua6�WW��voOQ��ÆD��pt�l
bP�&8�2}�EB���a6-n5N��9kiʊ7n���BF�p�G��B������3�w��K�I|��p�=���o�g]z��MHj"T���嫾�uՇ����� ��S�§��	Py��¸��n�g��	�*;~L�H6J�˻�Zע�����Jz0{/�wXk��&t"��%�ٓp��a����L�����8��`=W�jv]��ɑ��	mpa�.��$v3ΪD�����܉WƂ�*�&Jw�H�3��ã)$��3����Rq���1h�՘��'��dU]k�g�8��6{�؅I��٣ Af�%L@���Ѥ�f~�4)|�D�_p �w�E�Nt(g������*Cnb����6�Ek���\�w� 6ܗ%W|I)�&(�'r�K�N��7��Ņ����i��r���O6�H[}�I�̺�?��4�̕���cV	�% �\�����ѯ���b�Kt�����2"(Q)<�~�(9?m��D	�F���UX3��8�MNn����ʡ�"�)Ⳟ MѾ�(���ӂ�A���.�&@c/��[���Q�
}[ӕw����,����Y���}8��s!gB��?���H3�r�?S-{���C@pn��V��¹f�����ƪC���0��2E��Y睛�Z��Jݲ�˼�@����9��Pf��c-���/z��Y]"�|4$'b����W;�ͺ�]�K_�-�ɇDvPup��=T�л*|A��9=
;~`�X�O@�	�K��6c4����j�0&C�i��kդF�Uwא��9�jxh{t��D�8�!��GSy#ey�ݍi�_@���b�/*��EJjT��LJª�lo↨�5���ɗ�w�����9�>d����.�*�F0��0��j(LQ>)�ԥEc�'U�S�%t�-�
A�<�X2G��,R�ա��N�C�=a�`@��Xm���Gc�ļ��?��a8�f�H��K{e��r�̝k��W�G�{T��{I�I�%�=�J��������-���=R���h��
f�u����k�7֦���Xh��\�V=���ā�;�j�Yu{��'����� �ɯ�4�.��W�nh8D�e�Úo�'}�T�u`����&�&���*q~�E6��Vn^��.�&��9t,�7�,R�.�D�Ԧ��E����24 &���QiшKx�,�|it'������&��p�� >���7HkEb/*�SVau����vd� ��}Ů*Bq�W��22����bqt3)���م�a�P��Vw��)s���a[D,�Q���>r��-�w��5���b9��� Q�Mw��I)�أ�:]4<Q����VNc�)�Zϻ	�yښ�D�6�|�g�Z#��/��ĲD᳉;{fT�e�56��%�X��ˆ� *�P<� g��8������~JVWq�F�����
�N��iR����uB�nH���>m�G-�fo��e��1F���b��t��C�fѝ�B��"� ���������_�k_U_����B��V��ȡ	{�����4'�1qU�Ƃ��9��~����c���x<>�1��u�v4Y�O�tiHʜ�و�����w�^y�!����aܐH[��H	���LG���	a����Y�a߉׮�'h��?4��(|3ء^(s�f��3�dw�y�`D"���RPy*=9�IҦ�}?@r��\!i�����3��$
��k?��xşt�{w���1�\�ٓc�X�Y�ڑ�2(�3s�N^�O�`�ß�ѿ~/�;�Й�|����@� �J���G��nD
�Vdھ��&7%�����$
?4 *�<\��1,t��&�b�VTM���_��@����*8ܝ|���hm�>��oF����.%�il?w|��.��٭ ��a� J/�u�J`�-�Y}E�KF�g��h9��1��)!W�WE�V�gC�������T�0�)�ɑgҀN�?zc�y�Hnx�%��5?�j�~e��^Et۵=/kYO���?!����_�<�gF1q
�����|�P!Z��y���t���1ߎ��-m����3@�������N��.�l΅Zɂ�et��o��o<�6�t-�X��V�O�X)�,�F	��EY�2p��}r�b|� �Avލҹ�g٪a|���P�D���w����x �p9��a��^tX��^r�|P\[?�Fz�