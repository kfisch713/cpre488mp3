XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��K�9��z��,�Q5�h_ ��T1��`GN5+�Â�8b�Z�kܲ�nP]���"!}Wa���F��tᴲ>�V����Ҕ¿��k�������H��n��1b��N�y��zK�{����cj�~���~6X�8�3H�|�.�ZLψ@ъjeQrn�2⼪��܍)wT)e���h��y۪.A>�_>~�d� u�]�4?5�����I�Ppt�z��tv�C��.��sDWW*�A���T3$�ʄ�HlSČ����D��n�v�6E�HL�t��-Tbe �a����W��H��\�+5r��(#��S�T�+�k2�n����F�!^���Y{�>9�$2�8�i3���޴���i����Ei
�sh��3��� ��W�b�K{px��t�����q�rt�g�_-0���D��}~nn.���9���S�;S["2z�����J"�RH��C�k}�ŝ����t�򋡢���
��ߘ�C���K�&����tc��-�����*��!�iSG>s��Ƅ!�	�Y�Z72���͟��` ����#�I?������*2vN6�?�r�d���,�!�y�.D1��w5^O�#Zv�L~�e/;lcY��Fu���5n+c�p�XܹEZ�R6]���h�L3�T`̏p��B_w]�������X�wItM�~����D�������`z{��1	��m���s@R�`��f~~���ֽjh�ui���l�U����mw�6�h��WXlxVHYEB    3e93    10b0G<��I,�#�כ�e];H[�$��]��a��<~$�F1�<��Z�[�KO��y:N���!�ߜ�͌ژ�7�\�S}
�s���L���,�qo�^���l����8$�WOˋ�~y�ןu�x���ژ�;�(Me��r_��1�W��f���C����zR��=T����+�ϥ�.`>aF�I�5^���(���x���[��C�䬅-����*.�F\�l���U#�|��8��wS��U��&pn�`*@� �J���2��,��@&�F����" v���|��`	���P�ۊF�T�mSRpC�rL�S���~Ā�Q>a��R?�.[�e4�����g��I�����)��p�e��i�9��������sŅ >�' �@�3?\�D��z2cK�{~���:z-�����7��j�Q�O���DD�lgQ�W�l�����({",�Hā�K��!8��a� N�aM+>�*lٓ��y��D޺s-2{�\�1$��1������NW5��Eh]"��9�:-k��t\!�(k�"�^�u�ْ~5��!�BXC�>u?N!ZA`��y^j�VɰAd� ��2ɧD�0��^���{�@0��L�F��Lɩ~��-<�ոtPL�_��s7,x�O�}������{5�H���$)�=�J�S�[�9�!ɂM�k�2�)G�&���0Z#��"-���d��$��I��o��α��2�,F�]��e�WDa�v!���j�M����XP��2o�ev
��w�cfP%��Tt�;4�ݨ������ �07��!Nj._.�p�ʩ���S3_~����6h�фFi*��P�jT~s����u���RXCВ�R�m��G�p@
@l����(L��@��8*��{��z���>ʠ����|Ud�B�i�oH杶�=x�#��8���Na'�ݗ���}��&�U�ZQtY���'c|��
r#�%��̹15�;
k����2t4�e�r�r���֡��1�}�q.ˮ��������vn��6W�-���|=G]��Wa/���b~SG��:W/EKN�4&��)�6#Lkt��-��86s��*6r�s�RQ�j��&��U����]H;~��}��<�r3'"=(����O�D�(��:��Fx��$�3�A&~#�{K��u�̊y=�
��U�D�R]Ǹ�t�]&&��3�߳{�,�dT�C��yz��@��Zoʉ��׶Oڹ}/|ր��7���
�S�yF|-��YY�%���ޛ���T1�N�kGH�L��	�f51�p|X$�Y��i(�����z?�S�L>�[S��U 5��^�1��xU�vT�)B�J���N�Ef�lN� &�Ӭ���A�~�ƤQFl�g9[ ��R$�$��?����<4��|Q4�\�UDW|�$�;o��N3�t�t�&4��L՟�g�Â��t���ͳ�����<�f��n��B��c{^u�΍�Q?r$X�à��E�p�[z� ؗ�d�!f�I�×#��-Nr�y�<��n�1	����Y-�7�F�2�����(Y�mk9�e�)'bm�ɠe�<;l �v�J�vf~w��h���=^]��}Lo����l�Ţ�C��"�(��.�h�*�d��Æ�Ķf�5�Q�ZɊ,��w:n�����'��e����`W�m����㸲5}�J��Ү�'A_m���1�m{���W2�7�*Y�Р�m"�d���O�+�.�7�qo��E��0�28��O���OK��t �����B��wQ1ݔB���ˠ��>����1%ӽ�k�9B�!m�P��uq=C�� X�ً�@|^xWVO�.(���`����^� sZ�e���<iߪ�g��>�@~��%
���M�7T���EK5C�#�7X-B��*.��0"(��G�nPJ$�5�ۿ����SM����ֈ���$"�Z �L�� n�ɬ<bf�
�N7W��D����t���$����E�=�>z
>��=�0b*M1*evd^�q.�<�ީv��B@�6�t28��%�'�ß<��\�����b鿙�_&�D������ /y)E��P�~�ftۿr!��eŒ�q�
ȁO�l_��.��K����U�8"\�2�m��+a���(��^�i���b��듴\U�b�[ڄ4��Rٸl�_g���E�	U�����*\Bփ#Q�f>l��)r2�4��_�2�2��� �{�j����`��߮-�߁Q��"`본�||�����װ���d#�DɭK�����w��zA�2�`��$,�Vw�0�ϯ�����׷�n�#\�M\�3p��n����S��N�=���~PF�wf�Ã��V<b.�C�*�F��oӅ��CAf�l��σѵRj9?���䕬ӳ�|� �]�_$����4*����H4_�>�b�d��+���i�'��Y6/���V�-�����0��y��fa���WΦe'5<��%���=O��@ۄW�8��?����F�t��YU�5&uu�"x�2#�����jm����vbhjwaF��wD�UjZ���w�%YX5X(b�W}�䐟�N���8L:X�#2Ĉ��Y�U��"��jb�Y��7`Q�f�'��/=�mBo�0�^6o�n�=���W ޛ�R�E�u�"�'�z���U��%��H*Z���:3K;���^=)�r��l��[\0�T��zJ/�Dmֆ���O��%f�.c'��ݧ8��������:���r�'l�����c�SRMߪ4w:��Iy�ܶ@�?�<4X�Xʉf�`���\f:Y�g
I˩K��Z����+s$bV�Ii���7w���UR�Z��=ϵ��KJ��q�6��9n��xL�AÇ�X�a��DJ5���U�)�f�� 7�װ�K2oݖ��>�!h�E�qt��D�.��˭/������f�2bҁ��'4[����'K�ϑ�ɳ��A�9.�M�0��8~x���]�
)j�k��W E��|?_�,�Ayw�Va��?���|��^lCn���T��,K����5rˢU啖_����`�h7�4��@B��!��c�]�Y���ϰ�Mfv�՗���H���cb��� �=+~�D� ���<�bb�Dr��Q>�?�0Y ����189g�cL����c4�����U�Q����: k� pF)�o��Yx�I��B�ׄ����g�A����Ԣ0�R��ܔv��<�Ι���	�ʓN���w�U2���f:͉��ǥ*�H��|o�B�H/��d��E�B�l�X��C�y7cQ��m�}e(C9�S'�~(�^2���Q��*��{c0?�`[�_����'6���;:����8���:|���xE�H�h߁:-%�����/1�E� ���T��7a�9:��u��B[S�Q�e�
Ps��0�.�+���/]�����|y����'�a�N8>˂w���G"�L(��g�Ct���57��i򐸣�󥦶��/�������Pw������:���Ĥ8��D�Jk��H�� �@��4�s��Sǜī�pz뎐�H4>�0��|�6v��;"�inmW��M�e���6��V����
ͦWw��_4���D����i>�Zב�����܏�H�]*GS쳃�+��6�Kb����ˢ6��%Z* ��ݗq�`Ëb����]
��F�e�Fb8	�gG�̝�h:�ԵY��̬�`���|�Q��Nc��$�*���	K�\S��e\ÈbY	����su$Y�@�I��Z`*:!�no+דSft$F���K�q
{P��7%�ھ�B�u��an5;�^
�j��w ק��zS�0�
��G8�HN3Q4�t��HF�d5����RA���hݭ?��ϓ;���m?"�ow�ƂQF'�Y��/~�f����F���4i�kS�6�;���}}�f�iQ�znU����U��i
6T���J�f����N�_�LZ�ʺ���XTvP����_aPm��˵w�g)���xF��i��'2j�c��a0`}kYU,ӛ����!�����C8������K�#��A���t��������:�����;{��&��Z}��Q�^��ʋ�V �I�7���k68�q����L�g����52c����L�M-L|q<����-wW��sܷ���"V3V�y�(��$�� [�<�:G������3۟u%�Tܘ�v�)pe���![҈Ѥ�a