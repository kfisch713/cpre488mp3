XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�������< 6��߳�p'Y�ЌG�EkH�����ki����~��Z=s<~~�TU���^Z	�P��0��6��EiWǩ�J�aJ]��A?_鷎��9�}&���"�}@H��r]�h�Z3����Ӥ�Kg�$���%�����1Rkt�?���54IWp���a��Ġou~��K��t>���9���oWqa��&Z�����ק�Y��D�ٖk{cqUpr��w�8tĿ�\*����C�z����>�6(���9����kɟ�[1Z9��bܝ���֗�<ƍ�+��ݞ���Jȶ���;����µ����*�lx�v�qb���ۨ�߾���$O�̱�j	N�z�IBe�5��lp��?�j��e�~�q���M��,<�r�����|㢂
M��iyG�7��u����M�+zX�1�=,b�:�W�\y��(Bg�ׯ���kЯX�xi��S{��4���HJ�\����nZ�Wѐ,�Y�)m�Nx�Lf�n�FM��"��x���/���p!��a� o\@N�
{)�DX-\��9�iR�;�ϱ*OC7��@����N� ��B?�]��F�n�q�~b������Q��i
Ү�S�w�Y��nxkѷCg�Q���jP&L�"�̛���V�6�ͬZ��:��V�;���/�t�B�4�x��_K��o���?���9�N�����Ty.ZZ0�-�\���<`C��ܚ؞ 9p�'�Ma�pIQ}V�+J�Sv+�����=XlxVHYEB     f9d     6c0M��_F=�{d�|sG��)u�sI1e����{���8}�ҤLJ��#�wx-p�:iq��[���'�B	�$mľ,��Ճ����j�M��_RI�A(&!\aRˡ(}�lBf�KiVʹaJ/_RB/�DK�4J�0G�5!t�/��]�9Cr��%�ѣ�uR+"�J��A���t���0E�#1�W �bOܨٟ�d�D�I��:<��a4tGԖtP�$IR�ԏ�2_`���_��{E�������c<0޴Vpyo��>xx���n�������ED�<�f�܂��Z�9�����_������K��`�5|�l�(2��,wx��̸W�����c+��ř�m:i{RK�έ|��Pߔ���+?8:��XJz	�<.���R���6�JȍT����X�֥�(�Y+���o۸3��U��f$MM"&�]B�n�^E%�b��|���YԻ]�tP�ء3T?k!��`�:��?XR���˭��-m��m��]�H�6-�4��͟�_w,B6�1Fn�o �Zѳ�WD��Fr$惮ٞ-d��a��&��#@��5;��HVჰ�q]P��G>��>K�5)���a�S����,2�|�Y��I�>�7�8�c��GB��w�
q���P��P��k5܃�������nLB���u�2]|#F�Y��E� I��� ��f���ڿ^��a��EA� o���%��8���U�(~uv��p<�lZ��iV�jo�u��L4S��׋;J|�rW��{�6-�8��x�,_�!���&+&�<�zg ,�7(�P_��q�"tK1�
�6w�����r����քp����P[�`}�WO��:1�Z�M�CӇ[Ђ �-r��P���$S���|>��˞Ey�1
��G��qG�G����:��|	���y���
ԅ��$�A (��H���h�:~�[����[OL���4��!��	�.����`5���3\�K�``��iM��@�]�&�p�o��Ԣ� y���5��������~T��}�S�	 '�Ju���!�=|��_������N� ^��k��=�M���*�Ąi�T�z͙.Q��7ؠ�)�Tp!L��HoHy�(��(c:ߜ��@���;��-��4r�4�7��>�w���9�Q�OL5�*�u�ƈ�)����k�kC2�l����{�^�3?�����
�(PA�v�ݍ5�u�$��
���R���=Sߣ�F@4tT���:��L[
Dy%�%AGUh�	I���(t;��j��s&�wD��Z�n�� �Ό~樚��������=OF}l;�\� ǃ7�����jQ�aah'��Iڔ�%��,%�b~}Ͱ+���3|4���n`qa��׹�1�@�X�e��񑑿���G�^Ro�W	���8g�d�YET%�c�y�i�7��o{��k�K�$�޾�D�!\~�OBv���$U?�~�񏥟�CUv��j�zvo�>���R	V@?c��������?��B�K^�pŧS��x����
p|�s�4�x�6��v̢��9�3�k�`8�9�8��&3٨�]m�bO��*����?^��G��V���R|;���ɉ��0�����.��
p�?do�ʽ���O0O+�j�;nG
�"�T#T�$h�ҵ@��§�I=RN;�(w�<���{��c�}�z.���- 3U�>^��b�:�4