XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����	�6� �lY� _��W]�ս����͂�O,bc	Tf7��һ�,_�l-f�Ą:�ߴZM�D��s�����SW����mB?���f��C%��L��ܨ�� �*"%�w1�v�tp�%*/��xZdT^��`����-gX� A\�[�:������2!:��������8�N
�s_��<.M�7Rv��{Jug�U�����Æ ���R���\���g�t�ڝsJE/�7�~����#���j߁F~�"z���PgsiUy�O�:��8$���jK�c	
�S�|����FU�H !槓Cd�U>�^|ɠ!�	m�ھK��z�����;m%SQq8��4���|�ߵ�.�m�Ob�(��z4�`��������V���6W㙏z/�rY�+s({|��q�k
�c���Ԃe�ܕ|Wd��&��u�)g6����ޫ��+<�Y0<�����/S%c���uS�kjӃ�:]�[ mڈX'@Cg�J�Ӧ�!�9�
&i2�0Y?p��R���R���B��W�ʽ,!��D;�M��� ��j>�,[�6jD��Ttx�cw_�M�n�7U��0�*ƹ���k�D�����"�ے'�i�
������O�Rd��co&�#�D�c� 'Ŵ�#ע����hpS�p4t�h��r�[�K�u?�
0Z���;5�r�7���t3�����?1�����/
�Ԁٔ�?���X5L���09�ɽS$,{�.�����	XlxVHYEB    82c3    1970�t�t
Zpm�=K4,�1�=��Ѫ�_��G�a����K@���Ar�e��%h�r�mm�uEdPL@/��5�x�c+�T:!�6��LPS��-y@�]�C���k�]9�~��9^8g��ڹ����"߀wbY3 ���ɍ�E�fm�g��ǽSړB��(���q"��b��'?.����\y$�����Vw��BtB�- pX��k�������7A\���@�}h
Kz˺_V��{�Y\�TG�/�]�^ ��,���?����\lj�$6T��d���ʒ��A�.X�[q�/akb�ВA'�Y���^���=kc*�Rvl��!pAKIA-ia��ł�k��M�����HA��Q�(y9e�^�qb+ ��g�|!�N����T��ӊ?��ǫ�֔<���3'��Ǘ�g
��e}�-{�=x��A�����܌�G^F�E{ZZO�:]�DP7���3�p�Y����>�}��0APW�0����A��=�,ˉXx�C�@�}���%��q�Int��H�P�Y�(�U?�E�#>�Wp�t��iH�:a�v�5��:�]|��]�,�JR�dr�M1�*����\+����ƈ�vBɈ6��踆`���u�n׼1u�Ҙ�\ʨ���!��w��|+7���@D�ހ����D����n���	�p�:��4�K;�i�̮���ט`+�q����݊�u����In��2G;ZȆ	DZ�(.�3���+��s)���T�/�h����i$VL���s�?��\/�tA��.nF������獰��H~�N֦f��f/�P9F�~�n�}f�c���2�T
�VZ/�p�Rʥ���d���p�G�&�Zf����?xi����c����o�{�E�V�����~���"��(��������i����C���k̰���>�Rh����na�~iE6�=sT�R�]�U@:�O��><r2�Bl�->��Vm�u�ߩYo<���y���1������� P�ய;?�O�k�)��n��=�Q��
�Ä�(�i�R!��&Ϝ|A�u��sza@��.(!�7&��{��(�2�V�#��nx�̧-�c�O7�&�4Q�p��@t���֙�Ʃ�`�X<���=��P�����N3�Pr��2���h��(*�w���Uq���:��\ }�^ۇ�a����R�34C��3,72 �-��um8-X��iuzϰY2n�v0��<��������ۂ��xy@e�:�bo;�}�6�a�n�	1�!�,q-�T��n�[�РɪVz٠Gm�]շ+�4��WU�x7
��)����&���� �q;9����P�M�Rǔ��`�zr�;]ц#�P�������j�\X; 	��}�W�2�;ɱ���!0Y�#��SrdL'1K�2����R�A�B)CD�s����-�b����m��ڈ\�a^�-pn��?���s��JS��*G�o��Y��cY�Ă���;�ȝ���񢩈��mL�p�D�{ s*oSG����|�H�J����h+޴�X����2�\B�WO��Hs��59��j^R���'�4��H�N�``��ҋI� J��^��pk�Z��� ų��ęb�����L6�c�Uw���⦝�h���ć��E@zV�j������L�X�!HSɋ����� ~�g���O�����D��z���M8��DU�F/�S�4�hvn�p�D��\��Ƌr�aXD<�O\,����&�W
͇o��X���ӋW���҇D����W|�V��<-���=I�od���"<�7+�#��)s2k�W�t������\.p�5�	7�͌I=�Wg��Di�+)X�4���*{}�`Vs�?��8�X�8h=8q�5���}38��#"<�Ґ`��w��S.���W�H$�ϲ��9H�g�?��OX����8����!�� &�D?@[l1�纀��x�{Զv3VX�l����$�yq0b{.��g/+�nM�1Ft�/�ߔZ9�i/i;��Pݰf/qA�m,R����o�sf��A�X�D}��Zr_�� ��kh"�/�Q˵���=-��V%GѬ�Ew��%�#y9O��\����/���]��&i�c�D:f�{��{yWo����F�{q�r�U�����s�yLCR�7����,f^.4��f�;���Z5�z�N ���Lz=3ޯJ����t����ß��֨Ǳ,�`�g�-f���#1� �W%��y nXp�?��'�ǟN��}�	���L�.��(�4o�yej�UN_ۅ�`K1X�n�h7<���d��I��I�V��Ǆ7#0�`�^�E�"Q���$�ބ- ���7�u1>eAB+%yʳk)���;?e�d%��o�s���wfLP�wsno�,팒�֬�t�j����t0���ËL~y$������0M�6�F�m�/��JG��u�q@̜�I�����5
|���1w��KRA�͐}��`�+��r�i��ɂ,���	Ў3q�8dբ�퀧z�~WPS���0����flz��reM5^��ܦ&Aȓ���D�A���ᓊn��-��MWg�o��^��|6j`@��S�W�۾$�D#���q;����d������*��)8Bɤ�W�C��&�n;|[k"�t�d�ղ���8�&M�'��Mt��g�rvK��X�����z#��\�����b��/��:��[�(z�/��˖J���M�W�]�,f�m%M����}C,���֑����A�i�TF*yU����^5o��5vEL�U��Qh**�A�=vgM8[���j�i���GM{͖N9��m��kĪ��'�3���Nc���O��+�F1޼^J9zA��w+��~P]��Y����� [p��-��k�4�����S���ytZGT��<�yЂ_�D+�I"��T<�m}�[�"����,�H�G�Qpxܰ`�8Sl{��H>75��z��+c��g�*���e=�<������-���?w�?Җ��R�ԃ���z��a��\�a�wu,���0��A��W~C�j�� ��=��gճ\��jؽ���xK�S�AW�f� �JBC�G�TA��Κ��e�c= qv�s�k5Hg8��O�ٔ�|O��X��:<R;������`N����E#�-��`"*Ͱ�8��������-$D-f�-2��D����"t�j���Đ�������M��F���G�����B�5P���Rk�~�ȩ;hb*.�J-��:m���]��w��z��} ilܔ�ZY�0�hŰ���r�R�cw�/6]�� ���O�V�U���ej�-�dlQ%��o�uߋ�p�ᎆ� W2" 2`R9VEƹR��b�����ws�&�l�w*S���SY�������V��/1}���V(e%��(�
�������ʉR����䍃0�.  l'�v�}6"z��qf�Ŗ۲jǠ�]iS�,�tgB�>
�k�2Ӳ^��fw�����\e���]`3i��[6g{[A�	CӅy��s1�1�W��o+f��~�-s��	�JV�DO��������ka��v��pCz���b%�7'݂�����(��jZ���6���V�:���a2��{��ot4��3��	��k�M4��	�N�[Y�x�\v��
��;��s!F����-�\����ڢ&ݪ�a���כC� ڤ��	5D��k�d�ސaU:/x��q�Yw�]�rM��萡}zx���dt���0��Tk�B��H{}@�.m���>���$ib��T�d%��
F��l���U�׃Qe����3f�)~��q`$�s�A�D���w��[dY�v��1��㗊":2�p*xZF@L˓�����}��W�`�P6���? �[�ħό�L6�����@��w;M8�m�xl�&��KͶ*ܵ�Mh|��໩5�j�"/ތG�<@��c�EQD���C<ج��h��ʖ���je���>M�8�I�*1�3��-0��˪�J��]���F���N
�!�_	Tm��dt�t<� �"F�7/0V�2���8�`+�Fn��[Ec��_N����G���%�])1�����g����ƍ��W��Q򤃒�-���x����d+]y�יK��"Y��~�*q���P�d�=#*e�-:-�1��5/�Z]lE~���ւ(�
]��Y����Cd�K���ڴ��փ�-q��^=L@�����	�hK(8�m�Wp`eد9�ė+T����b��������o8�,�B�p���5E/���C	���`DB�WwCn��ui\PT�)�{X�zn��GDU�憬{���
�Qi!�����a������ā�e��O�&�� g3����/�(��ێ::$H)�k�n��#����sK?���\�:���"'��rߚl�U����BuD�7{Zo�w��³�& E�ǫQ�̔�X%M���ȺyF�������Ǻ>Y2戣B#0����Ӆ� x���N�Yx���Mw�Ǎ��vL�����ϔ��'��OzM����N8��Pc�a�ő�F��pA���F�ۈ�p	H)G8i�4p���4�ű�"�ǋ���t�0>*eKß��U�x̘�L�j��vQ�J��cA��<�Fu��F=:4*��ع�-D���:����!m��	R�I�˽u◵S�x#H�����;�Ȝ�Dg�F	K�fd;��#�}��Q�T����[�_~	T������pA�>��N�ugG-����D�XG�sҟ/M�C�l�v��:�W���[��*�55\�q�#5Ҿ�}�c�wv�=���5n�d�r�-���ɴ������lѧ����H��5$�\J�2v�5�P�S�O�d��hxT��Ft�p2n׳���5_��^�ƩrN#գ�<�鏟ύ����m��F)��4��(��)>g�{���Ǘf#e��ڹEH��]�
-O��R�۳�^C�/���_"	�	b�k��h�8��.U�~[2p��8�~���N���CW�k<¯��F�*+\�m��D;Q�z����"���yξ68���_F.�T?��*m�;[��CӦP�=��u��3���_.�c������HNW�A|v�=�	�UGR2�̩���q<��zOW�Y�N1�H��P[�}XQ�{Mb���K�s`b�.�6J��"�Ҙ;;x�3J��Bl��7Cr����H$��^n'ײ�[y���aw +@v} b�`����5b�98���
�[-�:AU����V���f�k��p�pu���E�u/��ݴ+�L�%��}�-�z��3W��G�fC_}h�fYtZD�
�B�6�o��=��y(t�4'(���/��ۄ8=X_�9�1z��>�/��Y����ˀAmR������G㽥:=�<�<Jx��x��Y�r���E0��T-�G�@r�'vP,z��CկiGؤ���`�WAn��g7�}!���z2���F����"0Ü�o����`���_8�9&�9�"�A�#���NK�Y<��·a�5��������j)�il;z�{@����ڦ넱M���p�bcI콴n&��vM�c�u�/e�� Ŝ��WC��K|}�~w�GF:�2����t�.N�;��Am�3�^k
Z � �Px��8m�HR��|�`��+��0b�����R
%�v�#�6ۊ��  9 ���[5Z�B��I�IYg
/�g��-<�[�|�Q.bKo�)�ƚ��d:���QQ����/)���<_!B -"���M�:�@W���ꍪ��FT���9��j�6���2�<ha�2��4}$Q"&�.d��qd������+<��p긳a��(u���co0ޗ�[2�Ab|#?��M�ǉ\���<rH4!�t x�kBh�ZuWZ�H_0�y�r���g)�Ղ�$hB%OQ4Y(5�I˛�'O��P;��;\5�'��i�E�<^�R<�z�\B>��hFz��0[�	VC��ھ���Ǝ�.��ai���ɧ�}i��؍U��t���^mxza�>�i �#z�v�,-SK�栜,�*�;��[ƿ���z�a�	��8%p����@fC�A�n�:��$�
��lHJ]�l���#�
?`�(]�j}�GEJ���>�S���ג��L�3�y�\�~�Ka�̦��8�`�@j=�o �+�~���Ia���x'abk���d3�}���,B�T���R��⊯F�Rw�:[V�I��C{�:�֣Xlc�Bo��\8����)� Kۃ�ͨJM���άC\����%���Qwj����ln�`>h�:��SCD���\����4���uų�e��<�bFn�Y�-͘=m/~�bxQ���+��u�͍BO$���$p�3���|�t��