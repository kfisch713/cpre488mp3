XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����] �;0HwL��@���?���0/��0��T,�US7j����f�C��O&��P5��5w�dk�L?2�Tă'�~������3�1���,pt��$�}�Y�+w�)���sF\��j  �������/�X�ٸ�e��h	ja������+֦�S�ֈ�#�=��f{_x$n��٩�SH����i�F���"�� ��54f@o~>m�;$s��*9�,t���̒}��Y��&��rf�u���V� 䟔�*9�VN�<<غ��0��)p?�(���Ӊ��6����ƫf�w`ZL
�D�D�<Ot�c�';� '�w{Xӊ�h:F2<D߲��3+���h&Z�ˤ��_X�YA���F�c��L��B?�+G�.�3!����8��s�6�V��?HA�טӖS't��S�Ӯ�iƿ�!����X�pL��N�:iq8a�ˆ�%y�f�\�!mĽ�ª���j�b玡���TL_��x}C�
T{�IpL�u�u����lB���K�j��������v7��/�aS���s���(�͡��IC`4ts�A�C{�d>�<'Q���ԧ$*ڐ��!�Fk��
������L�FB����́ũ��Ҁ=d
�R�
������dU�\:�f��K��Fg��k��*�/��S&&m7Z�CB�0Tsu�o$Ý��r�@������g"�{�ƀ|ur� 2��.k��E�j��ɽĻ]��J8!�!3�Ct+�=�T���B�s�(�4��"�0m�o�֤���PXlxVHYEB    aee7    1ab0�b���A����l�����cq�_>׷}�
���,�U�7��!#���CQ+ .�#�D(m7&�A;���y&�=�?���<=�ѥ�7[�܉4�O$�d�]����a���r !7R��� �;��/��	�0�.���ĉ{�1�vR6�%7�_�D�xs&+�_.\���z���f\IZ'3��9�H��ʎ�p��[��M��1ď�{/�3*P��Y'�����x8����6�`&�y���[6��i,Jo�@���̔*�X�"�#�V�J�l�˳]��H�i�O#�8�KA'���d�kj�a�-��#�t�x�
�]'&�z'�X��������o"|�~w�gd�oM�Ί���^Qw[�	^0?�%�.[˨�\(�nFNJ �KAgt}�=<zѴ�?�M$$p��|�q�o��]9�Y��6b���0I�1fgI��Z�nB7����������M�S�Z���S����aGK�p�~*-��Iq�l̐g�r���/�v�*�Ln����P�0��^>���R���Ő����)<9�<�Tި��UV)�J55��k["�U�>���}��(�ޏ�ښYMxPW�t2�-Ij}�9�;�1�&[�bt%��9ȇE�K�Dc��}��B�r�a5ꀑ^�k*�3Q����\c(�t{]��	��4$�a8xj��+`g���w^'�x��Iq�ed�{h�6
��ew�+I�s�jB�ٷ$�_�f��~�Ӧ��q�Pu�X�z�K�5�-ș�gi�q^�:Uc,=!c��x�bS�u�-
�bpc:J�ȍ,8��w��t�ߥX�H����Pn�cw��~+��(�F����=�u��?0[���X: 8� �ú;zĭ�J$�"�F�r6d�S���Ǟ���k���(�!X G��H�Tm"KS�Uyw��;�����Éy��-���_�2��&ԇ˙�t����4r�b�8��%�u1L�$~S�LklNk�
 �ג��������X�e�vޅ���	=Cε���!�N$��r�4т�b�3=��­%�q�Q��C����V�-փ�De�F (b�ηc21-f�Eg�����xqCMZ�ʞ.�>��-�̓�2�{�!C�6�bx��O��#� �xb��Ui��0�o�q�E�Gp�و��?�0 F��~�p�5.B	.�����L�<�s���x(�G#D��|,��އ��������d��ى�9S�F�p7��Xg;�8罌RXW���G]�Z�E��J!n�p��,_󗯍!�`T��z����-S?�^/��lQ��Կ>�0V�JD���L���^��]��]��ʪ+mʀ30<=a</��ߏnƵ}�����V��m�F���}F���9�ͶS�G	����N5h}�ܘ̓|I�͆#3��'�h:OM �BC�]<�0�C���� ��rDZҦ:�a�M�jUͿv�~r2��'��;���q���߶�y��Q�Mn�Z�pr괹ZM�I��hN��i9G���HM+�Md9��w�*����mb4PX�9�(�WZ+�k��ir/V\�Y���S�Ň�����p�²�}zm�P��돴�Q�H֛��=7pvK��9�y�U4��^ʕ����q9�d�2���rR�5�C������<� |�7+" �����|k���%���!d.2JO���95��v��ɖMɳs�r` �:+խ!m��v�P���^��G���QH5����6�4b��kK$tHK�A���{�.외!�J�K����}��N���	��m산l�������	G<�۞��Ϲw��F� E��	|�h�B��0.�E��3,�?%��fՌX��{��,8��R���ʑp��FVU��LKIg�����E얅�&��	�^�ް����{Z�&�臓�2'����~��e��� Wb=�y&8Xŝu������M�/;g�fMK`�v3-]�8������R����g�w��Һ�[�������S���ݠ�<�f����'���.״�ǈ�U�_�4��ϧl�%(�YpyR�d��wH_�C�i���/���/�gc�>3����0$&�*8�m#�����7����t���t�U�!:i�T����:3>4�Q=�ܺI������.G�mv��Q�G1�Ď��2O?�Ԡ���Ɣ���l��'R�/=Ǣ/����+��݀8*X�����!�F���5:�F�r�?��<��WqN�WA�N���z&z�r�T��&�Y��o��0o�CSl(�����{���ĝr�p��$��{S��$�3�"M��������M�,���-N7�5N��mΌ��?�s�M�P9DH��#FZ�\�-�}����Q+�yI�7 7y��,@3�! ��r�|�wc�)�
�_��NOc�@'Hwl�0.87C��*�z�JM�y�A>�N<_�k/��|�{�3�%�0�l�^ ~�=q}ն-�	�A���K�Z��l]޾И�V	���M1E!����U����ی��
�T�_��x찫���c�������x g5�(�D�$~_hU
���
�xl�׬��>��Q��4W(10�բ����Ĺ��=�Q�82��vF�Qy�ǰ�}�D���E~��֎:�F���̏�)o���26�L�<�|����s�8��Yj����W�΋5����f��jn3a�YO���$����a<����c�#(��������d"b��t�[>Hsf��@�?S��U\�%�]q���-`S��-��3F{`��~H�"��CJ�4�� �-�\�/p���nF�3����z�	� �yM���a!�мV �=@M�M��O6Ɔ��7��3�+�$�<����Z��2u.�u�Ƕ]����r8���fe5�C�<|�d�yf^���<~���C��3�^w�U@I:��t�>r� z8���:IV�w�䶧��>7��d�얨�RrH�^������ؘq_4.�d�4������X��U	o����r��>� +|x��p�ܝ�_W����M��t	��,x9���9|oB�衈�qB���q���Ӝ�@��1�0'{5�/�+u)�,��K`꩛Ϥp~\�^�0e���K3�{4���s�|�-��J�ȝ�t�0cы�Gʙ��n����4�C,V�<"��8FK�1��<I��39t��^"��`$���2�6��D<�Q2�"��b�^MpY�.��:��}���V���?,=��,�pl$/���v���L�|H'7+�Y����ߛd*���x���|��gW������#MI.���6E�oru���T!sb��`�^?�� �[�X���Qh��ɰ�-��
��:E?��	җ�UkՋH9�H*�e���KsIU����f=>�$RǼP4b��<�e��+AG{xwz�@ߠ#C�-�b�_��	�-�i�XvT;�O{�����}Z"in�� jW�|�~�2���h� �g���5/b���;�h2 �lb�p�1���C
�Q��{�n�������@B�&����3���KQ�Dܻ�dx!94��GG<� )��?Be]�K��Ϊ;k
�����k.醆��R��������6,�w�̈��e�^}��$�i뙂����#�[䮥,?/�a�E�`|���e\u�9WϺBi��k�U�#�.w�eU��ܚ{c�̃z�!8>I���]I�K�9;7����=�:=��S�#
`2�c�Q�I�1D�@NN4�Ps�( �Z=� )��7��h��s�$Ro;�+:�]��H4�:���G��Cu ��~į�5���n��C�q�^�S�0�f�CFj`?���E~Rw�]Z�
�T^�|���l�����;�7w����/�j�B����\�(Oa\�G����2U���! ��U��`h��B:m��eOP����gZhUK�O�I~#[��v~�s6����\�uܒ�{7VG�$�;C�}~���`A.y*K!�;N�ʞC��������Z��c�$�)��b\�@�a��da��I�k`B���yH�����몹�3Rb'jsZ	&�ϷU�/�ɞ�	"�UgO�<lL�����Ȁ�*�-]�`�D�(�7��$c �T-9��ӱt?Ҫ��J�j�u)��I�-/�&yQXi���cv�3C�ż
���'�:L�$�Ģ�\Z+�7�l�v���;"z(�M���	���ߕbr����>�v��@z�5�˴���襺W�B�Qs �"�(��Nt��κ������(<ݺ���x���(���n֣�K�L���[��&:���@A�;\����0�O�M�8���T���8Ȓ���oAn�/��Ɨ�h���a_6�f�%��W�Z���t�p��y��f�w:г��dٓU���%#T�]�#Op����#r���r1�W�HU��>��f~��>��KB���+Ҹ7H�-U��m�:bc�d�=��U�*/�֋J���-k��N��O��>�V�9i�>,sm�������F?L�_��ؙMi��U-���i�,�`;��B�@ň�9��G�+��FG_����``��[��1�8����e�R�۽�ۊ��蚼kb;@�Fj�bZ*)v;��M�{��,Py�ϫޑ���,�'�
�2�vA���b?��Ehg�a�cc� �yS;Ħ nr��g/��xO���?-�B������`��U������&�y��w/���x���t�&9���n�"�⤺���̤ii�T��Y�)�r=�.5!���F0�E� w?��Im\��VH�b����K�͍�*�6�𲎐U��q�:p>��5��6�hjߠ��]/Ǆ=`�	�k����1�d�K�BoH.4�s�1D-7�w,��CRb�n��XgD�|�j�sz��M����W˔�B'��X�+�K�r�Jj���V�y׎��������'�@C�7/vP���5�J�*�
�Xr�a�q�!�ȍ��`��B�E$�Q:�~�����Ǚ�)���q\ewȸm���DeVWs,���A*J&�Pں�hFx�B����=DN���d��#��^eA���L7k�p�j�NY��Iby޾��?�v�"����P`��]otka���ݦN��������	�PC+LB*�2)7��cSӛI���!mͼ��_/�.H��kQ7õy�>��ȕ�N@��8��h<*$m�r�||K�	��x:�u�8�]S���p���}�v�y��1	C_9��[�0��o�o���v�9������V7��.ye$wSlX#��0�c��AŨʼ��G�b@��e�,���Я/���E�����V�̾l[���ο^3�t�s����#�� ��?6]3Rz
�u�����ղߡH(2�?-�����
�B͘�b��T�~ɬ��Z�Y���gv4Ah��e���_���-�r#*U���5�ߖ���~)�}���N
ܧD�������
l��E 8&�$�H������n��n� �iU�9 /�[���t��V�Ն�n�=i|ܳ�q�iH�Y�!�-w�T֚sR`��14�vQ�4� /�am��N����/���x^����������-M�d�փ�m*�`�/:q���P���S��ͺ��
h(1�B���rqre��f�d>�Rؼ�
���Ӯ�	��w�.�ʖiM�j�i�3�v�,�B�<�#�bq��-l�ݺ������&���e%[�6rv�*����8{{�ϺǷ┡T�]�`6�H\�cɻ��&)R]�,�Ar?F'=��No���"�-B}e ?���g�"����SA����iJ{�e�ܤu�F`�G�����O�ds�`��i�ï����iI(4�""4���j���C"O�n�gs��(�K�c� �V���i��b�e^��%繋�Lʉx�s�8��]��
\�gY���r�/���?D����ؤH>������B�[2e΄~ҏ^��㫹���~�$Ev�J4W��=�XO������%c�|���;��`���H�A�Cj���ų�v�`<G���͠��l����ո�%*z���6E���Bk�C���_�Z���(9���Q��j-r>5�Q�	:���u�j�Ϫ�DWEQ=����f�	�>]�q�s��>�;�"��q���I�B� ���rkN|�Վ0�[���4�e˴>��Y.�+Ȅ�K�g��<�E,O�$;$%���Ҕ�x��B��Y/���������d۬*9*Q�-��C�Mi��w��H[�5���J�@nV��9c�]�l?��(�/f9����k	����KJ�Y�@ ��#Z�S꿨S�!`�^:�t���6��0z��s����]��|�]~p�9F��t��7��.�h��,9a�SX��fͦw�b�ߖ��J�!��2{� �[7������٘q���G����^FF���p����_�Z��7U`���(�9/��C��|o�
���Ho��qX�!�Y������"[R��f�$QD��ػ��<�8Ig�qC���.�i������8/H��tQ$�d,6�bڹ�xY�Lԥ�QC3���gU���������S9M(GV�Ѳ�뷇!��e���6�B��{��ά�.���5�ʽb���x��~uؕɩ�<�ő����eƀ�%�Ӄ_*u��h6+����8�YX��s��8�}�$�!�V�o����o]dr�������p��O�����׬�8^i���(�30)��j��o����[�l/���JE6J�3vA�9��X��l���>�!q[��t�D�p!�Z�:I�+�n�ܰ6A���܅g�X[P���