XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��v����7��=b�1�y�h��MF�L�sRY���
{����D�o_l��H�c���֙T�>:��?�OC�g��ٶo�f����}�_�yz}�8��v�������U�5�P�m���
,�����{W]��H""f����-|!����9�g'�F�v�n���d�A�;����Z�ҿ'���vWcԔ �b��8�JzI<��<bda1X �9"d�Ԟ8,@l��8�����쓍���֊�^�5������7�w(GY����~�	�7b-���Qv���s`~����p���8-���|����|��}z:�#����:+^E��w�
�����ߑ��@�1t��zp����/��|��}� .^��i��C��p���]5�� ��b-,��Pc�9#�QYW��h��T�Ƀ�P�'�*��q��m�:WL��ԏJޢ�i��N��O:��X3y<:/��hi��	q ��e�A�7e�LsMF�~�eX�&�������� {0�l�2�:{x��ECf]*�U>�'�c|���hv��	i�����;>���;�"0�b�fk�ȩ�y.e�8rF(�dj\�	�w0BfQ*���z��.\���ث�����^CKcC�lQ�W�W*r����32UE/��H�o��(��$�ϵkIWI�Ђ1��"<�n'X `� _.�,�l�J�1O��qZ�z�d�0�5�s�t�J	���$�'-����=�=XlxVHYEB    dd8f    2160��0��c��q���,t��.e�q$�bq���T{�M��H�U�}��'���F����vP$}|��?u~Qu�P6u�_ۆ2P�}������9�?�u�r�w�,�ǧ�g�$�*W� ?}�C򼊳$u���Z��$odz2�f�a�E��n�a�?K8ǫti�������}�KFA��:�K"[��O�ޕ���צ�?�{�<�{��G̽��Τ�<��j���w9�)�j~ad��?IX]�#���J��6q W4&�Y��şB��u��@�?9C���y����|vE40���	��GV�z�y>��{�)/�Ke\�<��ͷ�lLs��%[��'�?$kx?S��D����S�]��Սw��jH�49o�m�6m�0ɘ�(�\c��D�0��+����r0�8���?C4�=�����������&~5�l�#D��Y,��UHDR"i���T��4�w���u�)��P�GG鐔o�����b��aS�����i�����y-Ii��eC���vza����9�%���	:��%3]��s�@���ZgvW�s�����[>}xs��������2���rח��,��+�*�*�u�&%�w!7C�i�A�>���
_�z�tR~�ᆎ�+���b�8�c�׌F��J��I!�W��|Ǭ_�Ü���b��:R�sģ.uU�)��H"&hC=Gu���H��'��tF��:�����8N>�8Ͳ\@<���
У�5�.�r��_Kً����"�����&�c"����-I(i�D ���������z�#����u3�싎��r�{ J�2�td���ۀ7
�H�tI�A�'	�wH��O�K&��H W��- 9�а�s ��I�~��-���T\Q�������SO�wi�[�]Jb�*�e�Z��͸��Ǒ�\'q�`�%PҰ�Z2zGV5װ�q�9t�G)�:�$f� '����w�e���{v���WU�M�����N揶bn��=aF⻔ƽ?x�K����ce�_ҫ �҄l�%���X6굠�2\���L�Y���e�q��W�HQf�\$�K�4�Tf?�rXX�F�yG��9Ç��q^zl�0�#4U�>���_�I�/N�s
k�p�`sIkI��w��1����S�K��qe�
�}�1��Fq�����
#R�[C���|����,i0�p�U�X��R� [��.���p%�{���i��4��t��NI󗂔"��6�F�M�
���l���!2Y���H!"/<C�j{v|�M5#p�������U��. iD):A|��=�v٬�mxa{�U���GVO����+t볉�|c�o�:y3	���):CENT���~�/���kq?�S�%H����U�~>v�G\�C+�'t���ю�n�0!����Z�ә�@"�/��n��aјI���e�j�#w�2VM�K?,#ٴG�T1�7����2��?�۟W�S���o�Uយ��?z��mWvS�F��@�'e@k��]�_)�(+�:[h��ȳ��-�k��;�k�|Z6緢<�X&O��
�^+�!\3_�L�k�d\���૆?_Lٌ�����	7`HA�����J�t*���jo�M2���t0�``�w�,�u�ͮI+N(�zx��r��5ndt���CYŦw�/q�����t2�UXӽ�~T�☑-!y��z�v��}��I�1��w�!Eܐ�09�����\�H-eTt�2�c���e9e�-�Ȥ��3��N��l^\l�H�PO�|�H鞛�jNQ�A�R��8�3w�����?�^gp'���H��(���S��:�	LY�O��M�M�d�V>�^�����o�'�Q�A��^�r��D_w��L{����t R��X�vE�� d��G�b����PU�wi��eV28u�rpxv���L�K���8^q�ܚ��w���9�ROp�l���$鶊hE��Yj+�
:��`�L�,�'}�b�.{i����ٍ8�ƾ�#���
��֗�w�u�.zcRy�a�{�ݣW�X����K͘�V4��0>R�:[c�~[+��|wOV����H���X҄�GX�I���F������ p�g�d���}����'d���/�	�P1T;�K��W`KX����j��'�j?	�
/�D�ӳ)�5�D�'�+'䛮���5���rh�֤6�G*��d%�v�{�&s��rw=�������vֽcB��O@!�e�/p�y�N�����K�B�SW�|X`c=�-����'�
���"#�.׋�s<�#�GK^������e�#�������Qi��8���O�Ï��З �^?U��5�h�K@Ʉ��B��dV���Q�火heyǏ�R�0p.c� ��BW�f����lQ�O��
Fow-�6���"-U��䅦AQ�Ff|�p~!󦸖A�IB�b�85BW�m̢ b,ܧ[WN~�G�C��?��=��Mq�Al�l�
���E�k��,5,li���ИƊi��3p�,
0���㊶��߉n|Z��Un��t�}���,Ζ�������be�=�ٕy�!r�Iј���80	1�j�T0��Ŗ[�g�C�2�6T��7hYbwo`�zn�k&�۩��ң�!�)Kl���l��۔с�p�q�R͘ �#g�-�86�N���P�($D��e ���8[�3y��!H�3��6�XMR+3��)G����}��ŵ:�ۿ�+���&y�0�b?5�|���SAI������-^y������{Wb��ذ��GgNm�5Mhֳ��9���y�'�*�<^��+��l��5���9�}{bc�ԥݩq��}Q2����+��������#S9�p_rU����Y&�!���9�S�2^����ޡ	#̋��"[_?=��� ��ɚ��_M�)g`���W��Ri����ȼ�����x��O�1ǤËcZ���[zt����l<޷��fs�8ܫ yk���kK$⪺~]����U�{K��7\�p�\�� �7�O�/��c��>*��H�"˯E�TW�����{Ws�[��xX~��e��Z�sdoN_�$}���:�ٴ� �^�e���\l&�҂�� ���9'���0����J-{]y��H5���g:������Y��
Apҏ�Բd�*�)�`B���\1b�HٯF��E��"1�i%Y� :��Q)���cv�E�^��|��t���]7�9�Y|p6�\b�ʀ_I��s�]���M�4�Zꌸc�"�<#L��}��Y�/��,<���K�p_,C��N��4Á���LYҵO�#�(>��;I�ڨ�B���Gk���2�e�ώ;���籋T5K� �~BBh��0K��⽴�#�B6��r�	�/���+㚏��A0���i���#������[����ڐw'�4�����Zb�<z����yzwc�����qro��0�+���g���,�`Σ�H���*o���"��a�AǏ
:�b�!i�L��F֔�V蔫�Q�S��|#_8l��UE���^φ�|Q�ٵ{�����)T�,�'�H���8��Y��ZIY�SU'	������sw��ܟ?�=v���Q�~a�U��I�$�� ᜊ�g����M��<��%��!�+�FT,ħ���M;�V��m�S'I��U1V�ζ�-���y+�7
��,Z��:&u�+W��7u��HDN���m_��>�F|v���r�jr�oID�ta��m�:,qs�(a5��1 ZУQ{M��ɸ[M��[�#��S����s�By���V��^��e@��,&Y�֒������1b���+=�����ZjIp�.�<5_.��fi	��pbo���a��֨N��b�����\����q�����f\���_+��}]� m
U����r�Ȩ_�J��\'���,�&)\\�����a�����]��M��F����6���6h9Ӓg��,c����ţ��#yɧ0;��ZE]��UQ��t����V/�՜�������3Ѧ6�".�2���s��N����!�wnE��#����KYi�����J�u/���/�	�E�,�V�s岊�sI`�ȣ����gt?���9��O�[g9��u���k�s��p}�+#�cIʴ�8���|{fz�<j��ُp(;pi7&-����Ĥ�ۣ�,�'�#��`s W����3�švq�,Hr�����"Z,p�Z�?-�E��Ӹ�5O�Ka�$(-`s`TYz�cƓOO��$�K��J�ЋKOk0O��q�F�mE��8����Lw�Na� ��H~~�.�M�o	ь�|H����=;�B��Z��94����c�*?���gL�=m~��_�C��)d��c�6K�l'���$J���:�W���2�D�	��j5|�{��R�[\6bIyl���N<�	?���]��ڋ�b{�0��Q���3$���7fu��؊]��u�>}1���#��o���
�ڢ`��X9��#/Y��*f]���9r�绞���+����͓L�Ȋ~Uw)��i�m��t8e	��\3�T���]H��"b���*t��)<t�����h��$�BA��	�D�f��{y�Fa��O�R�m��h�i5k_6[} n\9�3-��.�T��Z��{��G�"_�"�����l`��ʪ���J
śM���v[g�(ﰭ@x��0)���,�34 z��NEc,ԝ2�"��'�Q�b��5�I�#?��D�����!�;v�cA�V��6D��WFqt%�t�yT�Ƣ�����pƻ0�P9�}8(���n�؍��c!2�Y������&�u�+����	G�gJ�H��YB�(�#�����*,%�L��F7�H�j���,�c��� ���MF��U��e4��lC����R��C�K[x�E)#��V3$UQp\mQ#)K������眅Rx�eէWM{���z�nqI�@_�����R}-@���������f�h�]�'te�s�g6�C�
�܍j#�ā��ӕ�-�o.A#�	��q����b�/@�E�!G1��I�PFa8ENy1��G{��B('���٢��&xf�Q����<siv8�+��/9v�"�#R*%rD�
�M~
�M�N��;��+Ƞ@�rN_��ۑ;�%Xy�G�.�k�4]�@b���quk�A"�TO�+DZr�����e$��6\2=�\Y����%�yǧدjĐf��P��"О�D��Ҫ�DOf}ЊwPv]׹"�p������2��	'����
)��H+�������L�'��`�.��6����T�?oYxޥ��ic��헇4��t�G��m�1 l%�)$ކz^�����n���E�Y�f]�ʋ�$�B���_&��{��71*�1�݁_��������r�f�@�{|���q;�qf'��J?��f�AE.F���'�bȤ�(b2�6�M-?�1bD�]���Ɠl��q;�oK!�ei�v�F;(����!x~Z=����\1H}�]CEdR�Bw�������Ǚ����]���*x�3av�*���������G���<���H��yy��oT�=�mU ��L��rg�J�'32`�r�"'?���FL�H>�G��9�e�
�p�]}Z���q�-M�d����\<1�r�O��>����nબ�Z��So����蚐��7�FQ�R)���:~Y1�r3ܸ����V!Ե�5⽒sR�y��ȱ�O�U��4;+p���}�D�E�GP��)C�ц�Y�x1�Q��)�q�L�}�@��R��г�G�~��w�z6����zD����L�'(}����B������U��b_��R>\������%�����r�n���DRR�����"��/Hv�B�yA.��Ċ���Y�o���_�0�0�k��q�gKes��,n��?��'NV��yD���2�fh�2�`!uԻ�ؽ�n0̔u�@s=Q.��2N��n��`�6������zC��6�����q�"�mK���,d�!��;U��q��@�ϩ�e9���M�>�
��alqx�#�#'z�=~�C�+�����'���t����KB�(G�0�*�4���3���j����!�+IҹNӡ�$��]+=+�3k��	]�3�t�;J����o>A���3��'~�p�䵂F��|����ǰ>�6<�����Z!�t�q��%��QN�0g���eQ�M��P�ݰ@(a��5R�y7X&K�V�6Ļ#<U7 �]�<�`��p��{���2�7-�Ca��'���b�m�����\ߵ�w����&� �,SOH� G}j�yƾ�I��!���#�dP�'����)��y��H13�N��u��Đ��8�X����:(1L�z��ե��R�ֻ��O�2�5�>��:QQO�w�^�Ԓ�'��y����h������?	?s4�1\		ZW��D0�����i' ]_�a��N�֊��~޵���R஺�L��v�x]^hA���� *��v�!C�I�@����NT8�_���[�G�!��r��5/h���s��L��W��-����+��Z�;�Ҍ�����#E�^A����/��&lG�X�/�Rv�/(Mo����f.�����O��=�� �.b�ʲ���#�e��e]�yV3�mRL*U�s���$ �T��(�E��Ri��r]�ao�#kw9��D�֖���/�@�J��fQ^���:���<�u=����V��[6�I���}`��LC_{�'�	e���n�!�w}�*d"�:�1zsU�O��ϸunɺ�%��^�2�Ȑд��o�[	�Whm>�������:��P4j.�:�����j���`�������Y6��T� �]P0/�$�&�R���=��Y��
]xQMºo�:�oX�%��H�u�����3i�!&�%�B�o�W��0��Z3#�s`��&�ѱ\7Ҳ��C����-"��i@h/�ɖC�R= vi�(����XG^��	̋����͢�\ƊAfw�yj���nfM
b�`��!�-�S{;��ʞ���`�c�&�@Sit�9���_�+<asځ���O�י^��:,�������{�^��|1J>���c�ʹp ��`� �;&��q6%�M�*���7�v�E)�����j�CS� >�� ���� ��؄VE�f���(����"ڐM���G������Z�Gioڼ0�����u��au5�ݷ�}�+>+лu��r�a���ڈ&#��>��	c��!���q7�:��X]:�]G+��S�):���-z.������[�� �"�`!+��Fv���4�����Z\C��������i�,�VAg�U������݊
o"Η�H�Ƈ�2��!�s�2����h�+Rp��@�P�J�@��`Zw.��bL2l�\3�H�ɳw��:K������Uw[T܂~T�Ǯ�qF{����A��Q	�'ت.ј8<������XX�a��V�����pyC���nIA�2���j�� ^:%�XX�w�(k��� vG�V\��4�4l��`��1l��?b�0�ʷ�&�:K��|$��w �*'*�	ۤ���˹��i{�E�Z��^���:z,/F���|�Or�;�pw�ά�e�9�E�/�I����h�FZw��(�C���(B���,�t{��Q� �]��Jcmp���x�@�0��A���O�߮C!��8e�9O�i���]����!Z3Ѱ���=v�#�˚��%C�'W�4�u�c�h:0��O����uE��N�t�A?"�dU���ΘX̵LX@��hi��L-�n��?����Y�Ͱ����]·���(��c�ڂ݇ސS?�=����M��Cؚ����Z��JXI�ϨA�T�*"��
���TL�r#��v�,LT�~S�C� \#	y�c���o��,���Z��aJ���qa��H�����}ԁĲ%�/ۖ��+z�v�w-j����B�{��e�FG�f|��#�	��=]��Q�?�2�0�t�ԍ��u�%�V�o�H�D9�Bm�(y���Ov����M�*�������#�dx�+sO*��(W�h��rȁ����,)2]*���(����9.�z�7@�4{ڜ�ג�Gr
h���P�T�B�x��T����{�J��Ȕ�<QmM@��;5�
锉�Ѯ��modoySf��v*�7�ʞ7��O������!Ɗ�����P�A���L�+ǖt|�j���M�i��`}^��u�k�~�	��=W`���%!�/$ې	LB6ۊi�z�6�J�n�|�~e2�Y�/6��)ہ��
�A��S�X}�Ԉ�^�Y��/���[�T%1�Rx������~�l�avDɍp{}��1�O�����_g@�Kzge��$��"`=M���<5���k{m