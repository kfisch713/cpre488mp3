XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�������t�J��f�����G��^��"��?��1�qKc�L��OEi_���0Q �Q��{���">v��Q�Er��)�}:�u����~�j��ҭ��t��QR�h!���]�����Ϡ�\�4��cr�� ��K��|q����I2f�4�ų�9b���� �+��7Ӗ�i[�yWqP�nT�V�Ț�a��6�6%m1��3�f2*��#�ΑS�p$�v�Qa��CC<b�cd�8
���V�h�H i��p��ɼ��	X��Zq:5�ٖ��Q������b���)!?�aᅮ�w{G��@��F�,��[��P��.]���!Ooaz;T�8��՝Xp�&`]�q����93��A�ckĚ��oi5�s�-�*p�A{U4J�> ��*gf����[�:���S�����:�c����(nx
U�g�,�p��R�&"����gV�o7��}��N[ C�;����mZG3����)���b�"V�{��֦���w�.��&K���ܝ^�h(��l���j�,͂�$;�y���S�v�� ��<8��d�x�]c Ɲ�H�:O�\���y��cB]���6�����Ux?뺴3Wϩ�W� "R D���{��K�F�.�.K�$O���Z��j�o���[reO�f1o�\�掮���
Iy���!b%V���MG�)
j��ه
>=��^sr�Qm��������i%��0�����I�i$�sSi��׼��ʱW�����1s�ވ�dL&���we; �XlxVHYEB    374e     ea0��ߟOxe8�%��e��v�l+r�QL)kk�ݲ�/�$Y@˱�% ~{�yӢ+�� ڝ��0ҌLY�!!z��H��mpCR6B3�Gf�@��E��PvQ�$������]�SUf��A����ň)C~K�')�C�w�IU�ݷ�I��
��.bh9ХɄE���2j-���xMUC�ţg�b���g7�b��w҉��z� �`�4��n9UARB䦼���C�^����*�?�n5��'5�"N���8V����Y����z9=��x��Z�!
�L�m�����D����V�:��X��$?�p�3�9�����L|3��w�#Ou���;�$�$m�����sMܙ���FA�u���Z6���׆#x��WYX�*�3D���If�Q!��=Ҷ���7��.Y����d���&- ����`2��fϩʲN�L8�(�m���F��WM�)Ռ��8U8Y�/9,��E_,����wZ�=OB�����@��cP�/����%��eނi_A�ivP SU����$����Z�h�lv��XZ�8�Gnk�s�.�4���8s�-�b=�f�1�w�&�`7�=r��0��iǜ~u��X�^����$�2ѨR��?����w�R��u��*�6�$c�#I�'��|%z
���jDuiZpVp�󥖜���)��:�VtF�B���Y��yK�����=�����^��fRh���P�7s\J�(��DN�O�~0-:�#B�mq����-D����N�V<����C�=�MA����m�cƝ�s7��H�"��Md���;B��x���v��x	�m��^�}�H&=OV@�c7X<���T�4�Wۘ�ݐd3a�3
�����H�,i2rG��Z�E7;@���N�6/�碭z�8�&j�u���oT�|x#W+��E���ks��]p=�2�D�h���:D��"V�s2�^�ό��E�����[_�%/����@�@�Y�b��!��&'���+�օ�l������R�e�`@�Q�+��/��L5ԥ�����^��g�6��k�Xd����>�C=Ij��KsOMy�"��H��6����f�4���D���0��}�Xmp�u?O�y�K��_��]U����S =݄[)>�_��Ԕ���O�	j$���Fοt��*!�mG�7�U���*$ˣ�9/�qg�="V,��ps�o�f\����3�8s�0�[��bf��N��f"���B�Z�
BE�M1����Q�1�����Y�x����Bѩ �$"FI���xB=b���dOu�R��{�t�� /D����LS��f,y>�wc���Q9��ⱱqځ�'5��
�d�'���̿���B{f��	8s�f8����t�h���s���M=	�ָ���T@iW�/�5�)E�a L��F��	QncI��ut����HDĊ�x�Pk9����b�"A�H���@��'�ź.�~cJ�0�e��8m�	 Y����T�w/G�Ւ�a�Ax��S[e�?��)Rl7�ǂR���}�k�-c�r�b������_��<<v���y{�k"M���c�Z~J�^�R�ą�L
@��1�-�Vmߌ�y�f5�'�K��^D����,��(Au�R/9z1Z�K*�[B�E�֋��9�f�2�W��U*�8NΖ�P˭~(��F�U���"�O�)C4w�s�` K���0~��@�W�?�M}����H�3��Y�vE:��l~�*>/�]p?Fl�*�M��<y/b~��R]�^6�b0Q@
� ��R�y����mBL����ԕv5E����C�']��-*�u[�l�մϜ�y��☣b'���!���#t�\[}ּ��O�n����并c�>���)I��3�/9q\e����^��\)V��y2,{�Pe&~_��3���H?����I�G#�s��(3?"��:��x�%>�T���~Ei
�?���,|�ܷ�Ӧ7,�z��O�?�@�م��YA���LB����3"VI4r�,��u[l�n��d�$֟��x�9��ٓ���K���uS�Ӟ��U�c���Q�h��D)t�����C�B���Sŧe'(I��:�Ƶc��>@4^�ˊ��Z>�͆��#�S��ۏ���*���_�k�����c(�����k�I�
�8���u�s�MlȊ4B�l�w���a��C�v��x`�O��O@w�.�"����`���|v�$��Jo��Ix�{�@e�C�?gծ!�-��|F�a�*}�5 �w�yz.��7q�Yv8�i`��L���� �����bD�1��n��� !�{�)����{�x����{<�R~�ñ��$����8�@./c��.�MȓK5�l�L�6M&!���*�{�N��Ŭ�\R+p, �U��l47�G�}�'��@����[��3����^��<-+�lv��n�K-*��j]����gK�%��3�N��Q/J���6 y�4�'՘��r�9�S+E�ڻn����ߛ���n&��;��p+Q�+��raCG��*d�|�E)-"	�5����} Nz�6�-l카�+?:ծP�k	9�0I�R=��hq[�0l/���j)� J�i���9:6~��E��%��.M"��� 	�b��W�R�z���Gr�4>�xE%�:����i����LN�@�_;�Ԫ��K��Ūr��u���=	�N&΅�Y�f�s����$�ba)� ]��<�������}�A��=G����P+f�H�������U�f�L¶�S8��N7a}��H��X�kp��] +m�P2x
}Gd���=�WeէnM)�c��O���{o!��k��×�H���9�B��Q1��8N[�����	�^Vf��U%?tlCXL�t�ʺv ��Z��{��ʼ�b��X�"$��%Ƽ�a{h�A�]y��Fz�A�GCw�C�iCicWq�7E��i�o����=bղ��*Q~ R��O[`;���ñ��\Cj�Qw���fV�)��ƃ�^U�.�����C�-��2wjx5���d4Yb����W��_�+.	0�_Ļ��q*���ȢW�
\207���p@� �0�L���l}����es����i�n�9rI��s��������}���x�b|��cv�P��9ӱ���'�kJ3�\���h�͑<��1��G-���qZ5��U:M�C�Y�*bb�$Զ�����a�R�R�t�w�������.�E==�s6��*{�Un�����岤�b]<�e���r���-� �~�Ȅ���a�[���}�Z��,;M�)�>Љ8����r�<�����ovm^t���""��v�:O��õ�W��5����aDh��㫽�$N?���Gx�$
�����`)y?�U*�"�����o�~=�@����F�1W�@y?���_9;&օ@�S����S�˗� ٢b6�哎w9I���hh{;Aͤ�]2��g��dlV�Eydx�P�d0�E�Q��#,�-Q9��x��Е���5h���߅w�v�Ǧ�fyI�r�_�t;�7]�IOA�0� �g�m�M$���'��賭|5��8�O�{��{7�E��XM��I�iU�6���hs`bФݤ�!��,��ǚ	�-��a?2�?8Ë�+ �I���Im�ا����?�R��#�B]���H��T����#�M~��TR�ך%�ӧr�