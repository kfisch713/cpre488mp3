XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ҳ`�������oj�{�.s�������8+Se;X:'W�Yj$ӎ��F������'4�����O8�z�=&\B���B]惐����yt�\�� vrq+Z��[7����v��'2���E����ks�>]Е��Iu!c=c^�����n�S�y.�i�AA��+/�����:NM��}�Xh_�dB�7&(��x�޴�;H@~َ,��C�>EZu�o�݅���Q��]Z��m�#d?T-'jN<>��3����9>�����瑶�0#dl�N���J�VS f(��� u!J�}��HqD}4�&/nU$e�z�86�_�h0��+�)'>�;6�(��ނ82*׎�aO������B��9�<���!r��.�q�]�s_�k��&7R�����y��r>Q�R+�A!� ��q�;`w��W�o �i��NZ)��^��0��� {�i�" {�ф5��胭{:��X�C�g���� ���t�FD�=����',�Ֆ�Y?���6^M�
�+C2z!B�P���R�OR�g�~v֝��o�e�7�"e���kBBY�{�������5nԐbql��t:�N�2��L[P�;pXX��D�m�q��2lҕ�� *��!1���v�pZ����N
t��[�>b\�<TL�M�#=٬'��c����eЗ����l�3����U{�Ԗ��m�К'��˱�	�n�bfv)Y+�)�\��Q���v��T��})l8uT�w>��Y�|�)�cw{XlxVHYEB    76a7    17c0o9�]���t�;Hӧ��̬]���xc�T�	|�)�́U8�=D8k�^������*����BR"%�n�L�6�d�#rנ��m}���G�I%O��2�R��3��:�+����5��j�7��
��4��;���X�|;�e����8��!pE �R�<3*c�)�n7M�0b�6>�羹}��͠��r������[e%��������� k�Ыqg�����)`��]�G���Y6�5o{1wb,��-{���R�S$a�^j��,8��l�oI�y1 :D�Q�hg�7�.�����귲Q|��rݑ��@����F��-�5�Q�63��&��ӎlǼG����a����{�Rn�Z�Z��.J#i�t�̖mv�M���s	B�:L�e'���GO�q*�d(3��W��	�Rb�tZ��`��û�wx �ִ !��:�� �m<.��|�����j�"=Fy�2J#�Q��]ݿu��R�������	 ~_�%�D����)([��7��tE�ZܟٚǰrN�t�^G
��'�A��bG��TS���?� ��yc��d�����&t�L�)Ҏ�G
���2�Au���^��<��G%�Ӊ�x^;��nZ�� p|����W~�'�Or2�\@W�F �t�,�AX���1��϶x0���3Ѣ�|�Le�;4P��$j^68ga�ԗ�oC_�	����2�9rЌ� �ձO�h�= �VEnH�/F�e`��J��4��Qw�/_,aY*�87�>Z虘��_��i�n8.���'-P�A;ق��k.z˞��*��?'�|?��2��UG��Q0J�aSZ���5�����N��m,0y"�d�ńE�w舘��J���	�ݶ�F?y��2�I/v)E�Ywɫ����2̜� ��C�:!A���W�;`>k`W�lG�]���sVi��V8���-RY�L�:�̢B�Z�,�:��	�`�ɩ�Gv�1�	34�7s�1��^�?����>6Әhr��rMО�7�J�4*�fJ��'j��;�veF���yJV� �<Lh�d�5��>iб@�n˃\y��Y���Ӣ�NUm_��7��3#�	"R�f��v���ɚ,2M��d�n="^���Z	\ދ2�?��+JNJ�����4^'�̕�Eq�W��Q7Fm�@d��N��Zh7@F�m!'
J*����e2}̀)�bj�m?	��r$e� �H��k����!�D`��I�\���͗���
O�ӁN#��aP���u��j^���<I���A�d�6��AD���� ��$<yIH,Y�q������A^���Ѡ�x��o���$�WƗz-NE���B�dR�5�$��V����lC�M⇡�æ6@�[�ˬJ�]DE��5`��L��9h/�#캂��}v��ő܃��.�-r3��c��4!�h`,�?`�
�٭G�+���S-�j���K�i�z��
*��i	1tW���y��x���]�Ź~���7pUx��y��z�:�Yh���R:8+�đǍČkї.ό�{�v�Ps�1)d�K�zf�>{�U�=|4�mVeחZ�?�]/,P7d4�L���f�w�{�
:�!� ���x!�o��eX�,���6����;�z.�W�%��d�Bc�?�Ss���ý�:��\_K�_���^���Ȼ~�]*����C9�㘻�SE��p;#�?���kO:Ҫ����j�v+-&�B~?�_�T:��N�* �Xo� �W�`�I����z��s3W2�+M��*����{|��ҥʄ}�\8�.�h�$yl����એȤ�=��ُ����׌��;�w������-��*y�{(g���N�]��[�1E�C��]'B�Ħ�,�B���r� }+)2jV(�u{�$r��0��Sӳ�`��H'?��Ջ�$W
EgD*H?>0���UK�0.@��>��)��f��9r�ӱ���a<_�T/c��}m�>2>�ރz�rݢ����<]�O�\��+$����Կ&1�s�r]���1&)��KX�m��u�k��%�ĠE��԰��y�{��n�3��L�;�'=�H�م��&14�9i}4
��ָjA�ZƂ��3�Fڸ(`|���:����V+��E���f�� tS�Z���rS*�Ɗ%6t��5�� ���������*�|[��'�;��i٤���F�5�)b�%65,�>w�v�Ǉ[�ү?Hӊ!�?|.���St !��.��wv� �"h�|�f��93���f-q�����1L�Y�D�L���$w!�+��7�c��X�t��;���_���w��rL��yn��d�StQAQwK}����B��9+\g�l���^�]A&��}ٛQ��V�8�)�Giŧ�#��|�%��HS��Oc��}:�QI����Hš)U��
#���لܚI��j�^��J*(ϧ_�Z;4��C\-�P|���Z~n/�����{���U��!��|�V��v�K��̞�RnD�o��D4y��9��fM~N��C�r��8�%Z]���/7�>㼃�dG�G���7��]��J�zz��ܩZ�q�C�B��ƵL�H䬕2����Aw�
�%#����m�kW��ȋ��.�k������"���ȏ�Y�/6�[$�� 
u�.������h�X��������"���1q���?�q�l��]8E�
�!|�g���l��Q���cB���cS<��^���֕\_�׆���P�W��@�V��]��3�\<�5Ce���fkt%s�|���⾉������t�V
0�:x1$��uނ��D*A.�ؕ���U��\1�v�.���o=��YT���<�cKG"4�g{*ɛ�K�� �������]�Q�XN(s6�%���}0�!vg��,����*d��g�s1�T����E�M"��h����ӣ��]�eE*�|��-' 6�R�i5�dO�1��rz��U��9<���(�\�c+�Bq�I"<� $$�l��)��Xn���޾������� 1�"f��6�����{�3�����$	�N��!�L����׿![\�s�2[ǷҢ&�B�r�]�	F3�Za�`���N�H��\��&�;LƲx�8��;����y���H��L��.٣���@��Z -��])T��Or�Vo_k�e�Ⰶw,z�
,xj���c��Ԧe_���sO�u��׏:�����I�������M;�v��|&�m�`��*����2PoM��o�({,�R�Hm'��Y�V�Ć��m��������@�*�e���7��i���Gfζ��Ď�{:Y�� gz6���G��f)
ӔP�mf^!�M��������2�K���>4��n3�[�N�Mc�殺��i��p犌����I"�����𚅒��!}�?�dW�ˢ
�X��*��i�O���!�"0dJ��ѷz�[�Р��8���87�*s$1׷ٻ�ӈ���=E�v��*Ӱ{[s!	n�f��a82�$N�V1�%آL,���=,1,����g�}�qJt�߽V���5��~���y�=�E�4eYݹ16L:6ג)�P�/�����~�Э��U����y����ys��1268�J����~,�"���b9X���ݶ��۵D�ų�8��g�ݾ1	�l��I�勛h\K����ր\�T�Q�/l%��T��o��T.��؎����ǝ|UnA�j��V+�"\���%�vRN�a�)���$6f��F/"V�&4���V���M+���[BƬ�.��D;P�3����ѫ>	�����Ҋ��d���V:�v_���uq ���[�*X�L�V����Kr�do«����u��[�"j���3��r���(H���WJZ�+�,�M��)������+=$�n`�g��������!}���/�{m�rN*wN(:���z��b�Ύ��%�.wf�+��"d�į'>{ר����Q)�����A������|���E��� ^~
t�qLY[��m���qN=��nD��{=1�CV�����\�?��}�a��H�Q�e��p8@	臥�Gb����h�X��-:ܪ{���a74�����ˀ�;v#�z/���K��W�y�.�b�eY�	�Eb��(�b"�1��yE['k�Fw�h���C��5:��Th��6M�b��}�ڪ'�a&R����z���t�@C���-k6t����-����8��ح �"T����Oߟ-j�8�G���e�^�j�P����-υ�vdf~��%�#)2MB�G��5M$��G����6�z9���am��U�A�A�eR9?�R��ǹ��_���:y��ϱ܎� |��hVΉnFϗ���b��p�/��B����M�����\n`�'�$���@ 0uB Z���~�YcB���k�X�2��]MM2{kࠔ4B	J�5�Y�<�g�5Q��D~UO�G"NW\+#��h����T�w��ؽ�M&�A�O�1k�z��49���p6� y�97�2�oW��@E���CDQ�ii�S7x"ϰ8<)[�"/��?�ᮦQČ�4D�g���uPz�r��GV��C2e|�|����@n0�$�x�0����u,+�D[>����
�}��-Ei+��4���2}>��%���u֤��#R��A�ep�ύe�:S~K3�u;��������Li��� ��K�z� ��^[���.ܬ���E�G���y�~
��K$�/T��bPa����V�n*׸�f ��Hf�G�Z��X-��f�oZp,��D�bp�鰂�a��49"r/K������0��L�`���� ��[��<�9y��`�vx�Q��ʥAQ��
rqo?�`y����<˾���o�r��	�@#����� d���f����^����^�㑕-�n���$&p���U�q��}ۊm��0;��:��"�?�!��3l�.��fq*�l�"��2�aZNk�>A�X��,(%��آ=����Ԯ[ZS�K	9�v�������3�,���g �<}9j�4��;�?�@~!J�^�p���Xx� ���6�6^�b/Z�5�ke)��\���ןq�6�pqD/X�j���V�c]��O30'�[�b� �t���_e%��Z�=;���c����f���գ(0ܧW�e�9����9�k_r��A��a�K6�M�x�h��R�L\�gI�c�/��Aզ�k��s�D��q#����r7����~�g��̕�x�4�kxT�8g�䥑�
�!N����᭭_�3!&���x��cuncd���i�6��el���j�_\"yn�a80���9�t�S�q	�Xh�偛t��c/+�R�8X����:ߗ2e�\�¾�Ǐ��1NT8�*勇)jJ������f^�f% /�pR�1 �ݑp1���:y}��г����{�d1$V �E�\�(�.���v�E��ή��zT��4oI�5
�M�0�:w�+��$�Ħ��9��(s%)���uS�����U�o�g��T�DD�9֧e�t�Έ�rΞ�����O/���'+tC�60_�،��H�D#)�L�m�L����s$D�W�o�׉��5�t�2�a�ʬ0(���8���K�<`O0��7����>bN\�ytR7~���ARsQP]Oy7/Q��"�1�ICN��Bl�Ns�D(Z����WYζ�G��WhV�<���l,�&�g�/Hᴆ��ךacwJrz��}���~�_2m(Ki>@.�C�j-e}�`��J+6#�w�nk� �N|Xm6y��{�v��5��ٗ�&��[�D���'X&�n	��+YA>7�AS��X̪�~zD�������{��ʴ��fG�w�&;*=b�`�9�K�|�!��?���S�����-�6����rq�a���u^����8�q�NO0�Oa��SO�=z���D��TVÌ
:��*��zx[o�2u.�n��s3���F/��"Г��[�Z���s