XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Ӟ#�$�\RCg�*6v�jb����ZxP�c����9��V}N�z�I��
�]��l� ZjG)�4��������	0ye�����Hί�-�*!,�e�� �`!�+Ta����*{$���c�M����:��y�V������H^;2g^A�mO�f/���As6����%��""�}O��x���^�Q�#��+ݐ�T��%Q��w�SkBG�	Pʉ��v������,�a��` y\Iȧ���^22��F��Y�7�$)��&�սFօ�U��v��縩#�s}c�W��mmTAU����5��)�����<��vQ�WZfw�v!x*� �C�CÝU\5�]O����M�g9���HUU�"���#���W�Q��(l����;	?��:_ic�ҬE+�>�gt>�\*�8\{A֦�n�=q�^ǆ��{���U���X/o�h��Ϧb�8v��5�~k��3��[�Z�Ma|�UJa9&���:��	P�t�%wq�'�S�S��Z2H�j��L��VKaL��+�l�C�f�q��|;`�*�q��������{��1��P}�d��ioI�w�@_#���t-IE��}���ǿ2$���
G��3z�N�h�Ws3Qef���긹
�44�����~��y�6�!��|�Y���'���3VkxЍڛ�*�ȼ��h���yR&{I�6ū�=���K�����M끏���-m�/��{�l�~��ݩ-����g\�刳���
�:�ꏲ�gh�XlxVHYEB    fa00    26e0D�e��ǝ�QGe+_�E��o��~X���߻)fzգ����	&}�8]��9G�c�@	��2*p����1��띅�����K)y��V�h:��4�a����Aю\}-�(�O���[V��n�����X�����A��֞a���P�A�r[8{!�}�z#��!���j�`�J��u�W��� �G��"J��0�go�d��� �Y||��9�GF��Μ;��������}��3�i�L��R��s�3z�3h(��)���2tc5��6|�����A#w_
�^�(����jN�\��'��1�d ���`�O��y� L
w�M����м�54���t!��Y�y%*��u�TZ:0�Z�ǰ�gn�+��P�G��۰Q�>W�љ��Z���H�ZD�Z�^l\�^~�X;�s�d:���ErT�Ø�$U޲�~e��c��6;>V�ZP5F���ݥ�M��J7Řۑo>i����x��Ь�%�+^^���I�����oi�΃5PK�(���|g�ަ����♨1Q���X�f�I�C���ǽ�90)�����x8��G�Ȼ��gdn�`H�f�hs��Y���ɱ~��l|'N��1���x�cvZ�uߖ�p����u�`2�`��+q_,�	{�6i�h��|�׎ �QQ&-�wVw�Kꆮ=(�(|e٪L-������k���{���8?F'0A�̅4I�dhM�$�T����ىlĻ�.�1m�����t��r��ϫ�7ILR�*pӡ���.��ެ|�����3��)��f=v�+h�����=�bR%�<��ɧ��xO����kY�N�CEA�Qg�7��/^�c�o�FI_��j5��`��������V��n�z��,�V;�Ȯ�4Mbv<Ŗ��^hdRh�������=� ����Ck�Bun?���4 �u�D�[7�X�F���b��C���1�g�@�x)��rG޵GX�+"-2�3�0sE�B����e?�.�&���=�ֲ�]Ь+H�T~�}��b��v�/��ԁ�I�$z����I�+۩�-
 ~W�U��/���Y��kg�P��=�v-�D��^�uׇ��R��rK����YnZ-��_w!��趖�6������0ъ$~���r�y���1�P��=�t ��^je)E!�wΧ�+iAdր��#���A�Eǻ�Ĭ�n��s�b�DR �_��!�`!�:��0���t���}`oV߾�)���P��+ �VD/Ri����D�ԔR���:غ2��N�)N~��((����N�a�qL�wi�[PB!e�E��(v����n�A��EX��n"��s�I3vp�øR�uz,Ua%�\�,U�4ScZ���E[y��y���_A�Wе���G�����E��MF܂���"�aQ��n�Pa {�>i*���d��$������ˁ��Ӧ��}���~�㧱j#-�1v�g?�a���<~}�G��KA�=��0j���w�([�I�54=.X"��_�^LQ5��0��5�M�*@ϥ)���A��§6���O9�?��O��X�
ɶ6Q$�˺�|J;,{�����u�x��0O���݅�Hf5}|)�>�H��怳�Ȏ(�!;�Qy�������4ئ���	SVT6\��C��D���4���>Q2�q��8��3�-Ɗ�'�	
�hM,Ŗۛ)�'7��˽u� ]~��'0��{�U5�9���{x/<$Y��j��~(�E��\#uP�i��_�4Y�
�%}tn�8vj����|�=����7ч�_�9R5�{�vO����M_ci�5_�L��gG�qg�y��Kħ6#�1��O��~��E=��Ph�c�'�6x]2؈�����MG���1d#�/��m�u���*t!���?AE�쭅R@�������[n�+%
�Vۍ�ա�Z��D)�9O�hep2i@���~���;{����HNZp�!P��A���-�ȫ\�3D��Ƀ��_�V@���"{(���&�f��K&�٧�iJt9lݾS�6�U��&����9$�&�����9�����O���	���Q���cc�,?k�@�S�-0ց�҉�X�~ǌ|�㖓������E�=�L��8�bK��!��i#�҂��mX�)��de�^O��j1�NN�suC>�)tK��?� �V!5j�*����*�抲Y�[��۱�钸d�U�?;.�>B��Tv�{�EWN�ע�Ue܃3*� _+�=��:�yDϽ���#�E,����"�rp�����qG��L�v
�?�v����W��?~�[�AV#]�=D�ߣ	�]�gDrM;D��&݇Y�=P_��,��xe9=#c��q�JI�y��ߺ��I29���V�����F+�h����#r�0���D�O��Ѕ��W[���� ;ICl�Ήŏ������_��Z���i7&��%�w�IJ25�T��0TS	��X�O(�g���d�,oi�����Kiy��/�����p(nO$���ܟ�2�!WKs�o��I�7�z��e�L��+���u*�LH8m�3�6�i[nM�])��Hϻ���-�����3����d/k�P�̯�2��]p���N�YESB�	�d�x��qL������UhY�2^/�fs���yҐ�������]���^�*�hQZ��W�ko���D�N9@�~@]��FP��j��O1�X���[����G�pt�$��t��*~5��E������m?��!�Ĕ���UF Z.�����z���-K~>�C����s��f�R�Jh���n���o����$Kk�_��WJJ��O
p�m[�4�a�d��>
J��K�g�-q|�?�m���$^�y)�R^�dna�h��\��
X�sOth\�V�^r�q%�Qr��e˚zб[��<;����_�Wq�-�Q���S�B�X< �vӻ��$׬��?W�>�On�Yd{.���q�֠����osv)������;���WJN}��YB<52��ˋ\��PW�f]�(�|<�T7��FX��e�hM��l+�� �h�	t�����[�h;/c���xxiʓj�.��
���d�	|S����qC��i2{4���J)�E�Y,�	�5��k�^)��Y�)�(�N</���BM��K<�)�XS�`&ã��Y4ƈ+�� Sv���m�*M�di��=���-�>:e��fG��1�E�n����l�2	.v6�_g��U㯢t�p"\�3s~��wF({~k%�J��7�_L����c�.x[����"�D�hj�n�p�:{Y��H��������F��V��t.� D��;ڌb&���y�|�k+1t���89�r��&�A����I�y8����̩9J��/�@8�Ćn�Nw�,��ĝ����=5LK3\�n�"p!�Xuw��j�[<P}c�]�#�wt<��fN���&KVl�n/v���@��lj�s�!�R���ł=�ܖ^+�h����Eҧ2CNG��l~�)�&���;"a8�����6��q�����9�"�.�`�zI�uTȳ#��=&��B�Ύ6FM_���ɮ~����?~q�����Ӽ:9b4B$�C�~���:�\+^|=��Mݤ�����ڨ������]/�ԛ���g.+O���G�Mt�F���aE�x��T�%L���=�s3QE�>�h��r�0q�<�d:�no:�>\����_oҤ��@�S��[M7�O�)	���5ĸ�S7��'�w��_��?�%«��S��W�?ᶫ#a�  ��lwX�?��K�(?׽��ǋ�*�F-w�!P�"�Ƴ���H<e:����x�VK�����R�D ���ч�='��:�qCOŴ,��63����p���#�0�^���4?���f�l8/�0�X�g�7��p�7�j�j()�t#����ZhF�1�[ħ��g�L�����\�礃a@S�d�|�)vkQ2�u���B���A�+qfo�%���L��(� m����g;/NG��Z���R�j����������v��+����W�v�U�9C�̘�m-����S�(�;� dL�=d_����kO�y��bR�V3J��i��u���1�f�!|z4��d%2e���tǄ����\z��=���&9=��ʅb�;>�JZHLŉ�Y����h7�	-a�;Uk��?h�e�`�k��\H�t��xƀŝ�}��}�X1�<ٟ��bUD���p]J���i_׭m��.�v�Y-�S�����`!ؤF�b�ٲ����\�lxv*�ᒒ���(�%���^1���7���#�?6@�-z��N�[��>� �����N������]7�
I8GA�٪ u�c�9ҕ6*�%H�{7��]k��Ȉq�z,������iL�:�����2�hL!k?kC��s9�6��X3�2�,����B��t$> b��ʞ�T�b�A��Z��$BPNE~Tlѱ"�6�S�c��e�Q���7^^�����%�2$��ȑ��:f�l<d��w��9����P��]C}O���វ	H�x�`�ƴ.Wl/)�@	b�D����$M[2�[� ��R��Mٓ�3����K�{��ӃW��x����Q��iؿv�2����0(���(�0y���@F��_[���T�nPF0^���=#B��V�v]0^�s��is�}��uۖ�d�h�9��7�"-q�,(|]8����'�{��J��+��/!U��-�{��h �)[��l-w�����s��rm�=H�:��}`('�q��v5Y�]-�U�"9߆n�����%����{~�dfwg>1k��	jom��)6�&�� ����2^�W�Ԟ���&a�Cz�^s8�L�$��Bn�%E�ʟu�R�9��\��50r3?%�/�|W2?u�<��T�>�BYz����zo���H�h��&a��[t"6�ӊYC��C�LnD�)D��tm�`��x.�35��4�2��]�j���W����Yo�6b�,樱!&P�)�� �6��ڋ��Fꏢ���j���E,z�u3��r [[�8X�,�m2ٙh�q&��:>���o/��y.�IVrr	.t2{j��@�w���Y+����HM�2a.�B_�Iae���e3�� e��	}Qu.7��KefHn�ڹ����ϘFI��r/�qk��'_�s��Vn�찕,�L�Gk��.`�=ε2�w��c�Å�]�q#.�TGA�&���8�u.\�������!ؘ��W����&		���;zs\�V���{|^�R����璗MB�ye�x�>�N3���%*��m@ou+RI,�6WWO���$�B"N�$O#;�'�B�m���O* #lN�=����F�1ڇW�����1��0�����)�=�>{�*�2�G�v��_t�Dj�N N=��&n|����КI�̒�4S.T>��"࿗iީv�g�� ��v���N"B�d�à���Ҽmo��-���R����G҄��B��{��{7��gӁq��4����G��r9�@{�u���PX5{��;:�|��mG��#Tza"���h��"��ڊ���-��[��L�ߨ������I��o��q�Ldb�e"O�j�V"���(�@s��bRp5�%��_�¹U6fws����]���{�vI�v<�#+t~[�=���U�*�F���k�hb��#���X�(G�<
�C��>iA+ަ>䳪��u����&G�kl��3��g}L�U��2���Wq(�ư��c����X�@�C�cbAĝ�TX���qovl�y����ڕͻ�q��O����Zݽ�9݋���ej$eU���S���!d�#�ʶ�]��h�AVx��i�'&��;�y����n!^}WV���;5֞s�Pk��L�TT�JB��Σ�Ђ�.��'C!LXFGy\�}tV��[~��O띩ߓaY��=��7���?��yT�� ���l\��U�� �մ׫C�����&:ζt���#o�|���0�9�I�ӣ��y���I��ZG�8������9��4U3����I���K�V-��i�P'�_����r����`;���6&|h��k����9�Y`*9��$b�T1�,oO>�z4�+��#�?��eu�"�.[��,�n�G�h�8�����ѵ)W�P���봐�(Yc��^���U����W*)i�ʔ�\�`C��J�*����^�����Gv|m�џX#�����+P3χ쐮qR���=Ԃ��L�����ƋЁ�+1���@ɾ�{=��tT�;�,�Zp!���p�1P6�H��+}�y>��ء���OJs�L1��g�\���[Be$q8$���8`M�GWF�#�\t\i���`�*��ŷ7@~0W��Pi������g	�i�	�xf�.�u��vKo8!�T���}��nu����r�Hi��i��G��g�p���p�R��i^���P�
	s�;�)�N��M�L��Uq��B2�s�$�>����)�Cu=N���Nb�!H+�?;�^�/��H���ל&D4H_쉛�I�-�*�G�1�W���F�WȤ�:4_�Ph�ۜ%�~�N�K^��F��b7w��x����V���Z`Tܿ��Z6 �OE=��m�W�!j�7t�s�`��^����@+������.�|?���*p�+9�o:x��-��=[>ZF�z����)�����nЏ��qǝ�55ز<c�l��D���-0Ўa
L��J�>�^�dύ�Iq1��{]p�C�F��W�����2q�ki��`e�1��HԶ=����6�6��ͽ�d܊��fP:!�q:6,v��TfB��|GG�u(�F�{re����%38`��E5k�y(�z5ګ�E��Uk���z�G���+�?p���DNark9 ���3��c��Bl���wM aq����	RgK �K;��L}D`��i��.��ak�	I�h�|�
�o���Z��塬��휑�&�k� Z�������R߈�D%_�P�Mj����t/ч/�y e�������&LHhK�
�}�Sͺ��["|f,u��~�^IM�~�&��>��CI�!�9D�T���M��L�����d����3jxTzd�8%��tѶ���/����b[��(�z�@��}F�[h'i��|
WTA���Pn-�w���'�ɋIqCʆ�.Y�a��h�z�Bd���;��@�ē�ɬ+}�w'��O��c������Aad:K�L���e�)�R�)F^���;`���_l,��ƺvpB�X�#1����
^}�����������Q:�4tt��,{���ד"������~"�&�pg�Mz9���P��'J�u���nmP��� ��R��H��%�6,g?~�Ej�$0D�4P�qj .��Ss�4)�� �Ӛ�?ꎾ9��{�Є�/����I�L���V��pO�ܨ��
d��3�~�~�h�2��v��"���P��zp��
2�g9n�qA�,�EA�z�\w�n��7=��T�Q���!�}]Y4s�8u�U�U�Z���H&0,E�8>ġȤ?�
&5A�0ٔ]Li؛�Y�����Wg���wVsgZ��ĕb�������v���N8���V�YB��R.��L�A^��B����-����S5kW
�<�|���|扗VW�������=�j�*�ĭ�=���@A��g��4?�֤7��n��<�fu7�2E�W>�W���!�K�#��mgMɧ�� �.�W{{iz��3�K�6���߈v��CIءY�`��Ak3�~2�f��HI�	r6�d��P��@*������U��cǙ�����7���_�vaӾ
��s��q��|�\ݥ�.�T��X2魹��lsYT͠��@�I�εX*���+{��5��ߐTM�ʠ���D����֨�����;�E���2I�g�efc&a�Ģ�#q��0��j���~���1^3b�%?��u�i~��ލ�Ҵ�r2��@`���.��{.�a-����́4sf_'�앞��\^���
�-1Q>�������\�>ȏAG������T>l���_�9�$2`���l�;9�T=�'��-�C\�3��g*��,�/=m�����ZF���Z4�o���O����RR`��wQ4^n/�j�7����2��;�����7Gv���X�_���6�t�O��r�0�X �m��Jv�B�⟍��ᶍ5�;��>g�>�Z"��Qf@�(��Է)�e�!�൥����^6��G~�Dg�!��d�0ي��?nMEY�3`��>�1O�~�8n�;�Nn��\6��l���s6��(H�\K^�|O��Z2��)��p���o��{W��UةXI��s�ŝ��q�En��J,�>���7!��猏� |�9��v��4��ȶ�6Ni�D� ��=�
�����oj�.�ލ�H�_�N�̮�I�_ lǯ�ʙU�%k��1vJ.<@��"K�L�+~i�ӹ��dʚ|#5&0�����hP��F�\V*�c���Ap�������D˷Y��4���{9i�B�$X�]��Z��(2tqv#c���NI���X���%�0��P��LV���M2�b�3C�1o��l߳�=o!T��"e7��Qϻ;A�,�D#�t�4�|RE��XbE5�|�������P��*�	�#]ʜ���?�ń'-`��i����3,a{=��x�Ό��6��:>�LF^��R=D>u~
Er�:@�/�K��������.�k�zX)>6}\y�nj��^��"�o0r��,>��X���s6���$�������T1�K8������4/�ԥ�ۢv�1��?��%�%WoE�ŔC8�<=����C��� <�<p�z�GřZ�$	�F��t�&_��:�L�R�G��ޠ'R�)��_[4g:Vs;!��LuR9)����>m9p�^�XA�*l��{��!Z� �5���?�ɰzB,UWi�?W���?V����)�u\κ�&��u9���6Mu����w�
*tY�3�>`R�� ��̝l�+�Dh���:}�_x�����E��8
#\���� �z�<D������<��g�H��C��F�G����(r_	#"X�~���{�@���� �����m=di��l��;Y���VbW��mQ�nf�������7�n^�A!w��V��]��X�t���26X�2��ح��t�;Q�4�v���q��l� ׎�_�I� qȳQ/�z'`$bH5����%@c����gbA(6鈗n?�s��ߐ�>�N���ת�co�s��>OHv�ݯo�\/����[��S�������<κV�{"���چ�Gm��!pM@ �X�g�I��K�X�B^JB�ˋ����vO����Q˧���-;\G���)�"n���(EKS�|HD�c����t��k� �W�a\m%�Ц�i�?�h�b�u\9A�/Qe��n� .܄���s�\��A-R�$'l4!� ��#���5�(�����ą]��*[�3d�8`Pv�)����7	����-���m|3�������+K�M0}6�,�����9s�\ԉ��K*����9T��@X��q��9�,��J��A:K�  ͷh��F8����V� /��Q��O���.;DԹ
FwA�Z�g��עʊ��/T��ʗܳ%�+h�J��
n1\Gc�/��M�� O̲�К^Z?����"m��bngƝ(���Sv^tӯ�#�I���� `���h�w��F���4��K��5T|� ���y/��)^c<�@�Z9xN� ������df�����F���Q5��{v9�i��Qm�זZ��H���MfXlxVHYEB    7d55    1450�bF
9�F���w�0��ԆE~��BN�Z�#YD�yj�q�ʓ6��J�T�������6.L�Q����w�i�y�����-i�Q�1���Z���Ip���J����I�']�Y�0�ֺ�j:�o	5x��C}aW��Ls��`r�7.�C5L��ߙ���U��D���:�z,��?�@d��w��ɇO.�O�'O��$f�7)�H��׫��N��ܫ�i��p��]/��2��&>��������{H��:�3�3V�w�J#.T/��dv[a�Eݎ閱3! ��ׅN:0������ƒM� ~�����{P�ׅ��0�����x;���c�S�-��T���/�϶��dzO�.MX?h:�v�W��L�̮X�(}���P���N����#�כ�c����xl�����d�Y=�wf�#���U���k�9�	Vn�Y��T���%�r��HU���0n�,����]0Ç����-üT�F�$yxfs����Wh��L������ᶐ��]^��y�F��T�p���(�7ɧ2Э�J�dh-�=?�'���/�$�l��s@���~����3������"�����U�<8�J�8���[����gԧ�&TX&��7N}=l�7'�!�Q��{5Q��J�8�p9 qw!�{�q�,{m�F�u���U���a��� �S�q#�'�X�ӵ,¡�8��]�P.�=�JI�Q��O���?��QE��;�a��c=�;���ak�\� ,����Vyù|�ul�+�h���	�~o�:L+�T$]60�oꈼo``h.�` ��ol�����p�� |(�S�41�k:�S'Q)]�&�:O��o`訆��}d۶��m�(S�WA������n�R qYA`NN��P$�a	Dڰ9A��y��b� "	���ڶU��͑�1{[CP��ȇ �X��u�����Mt� �<�P������\{����PnԻ�a1��h�,O|Ʈ���`�	@�5ֲ�ۚ��A��S�Ҷt����2cج��d�#�5+����P��0��?:{���~6m&+Z���J2��;��{I����A�~s42��%�Y�Աr�4n��ܗQ�5"$)'b^�(������F�r��|yH�/�>�@�� #I�C%ag�밾-�����B��g�Թ�H�e�-��Y� u��K�Śt�������6�K'ո]13�,�*|�q�
�x��1�����dT{ُI]*��V����2t�>�b͵�3BTݹbl�:�:���4k���X��)��g�;�ţG���͗�7d���gBV���!�0���<6����a1������}�{�����Qi�m�qx�.�����-
H�4�zO�sR��Ȗ���;RZ��	QaS�[$x�녖�_\��/+3�A���o6���X��z	���i7��^>η�G�	�V�=b4|1	H9
m���\�Kp�5��Yd�^�M�����?*����m9WF�1x饭2�,�.&V"=�@`ͣz�������(s�d���[���\i3�A��,`��AГU.=�>�iʛ(�ײ���&	�p�mSf�<v�c��%^���a�-���Ҕ��F\ԅ����תT}�7m8hF�0{®��J���sٕ~��d�����wx!�w��N�i�a�Q�����3dsf�N�G�1�>,��D+��+"�ưjuW�Jwa��	��ǛLE>
Wh߉��[�M�=��2^�o��I�,D����E��AB�z��S����֭X`G"u��������j�Y����Nc/Sv��A'
�H~A��&�w�;��mr'{�8
PŪ��`�X.�I	JI��4\G�mO#��re���JK-WWp�4c���0p�)�Z�X!+�P<�_������i�X9�
��P�Z7�%��ۻ���7	f�z��ڧf��� ���-ze�Ä��s `b� �P��-#,�j J��m������!Jh�#Oђy�ɍY
��ql�d;?�zK��dq�R����_g^w~׽�p�����"y6���cIR&�����hv��h1�	;z'����]2�	մ�)�&���D���~4�k]֕ �[YU��b�f��QB��d�HߞP�k�_SY��b�sѡ@`H�}���W���x�E�?�����S��l��,,��D�m�K��]��
���g�D��0G��J��k�A:z��,v�kd��o�'B*������6١�e�(eC]o\��)��w�'�W���K��`� �Yx��n��!��v�Oܐ��?:�
u����;F46�y�ۏro\Y�A�a*3` 1���>���!��Fb�3 Oh�f�F����OFQw�B���|I?u[�6T���������CW6��_M�%��F:ɇ��n�>��O�����^�I�I���&m���T{�>��Z	�;��ԫֵ���j˨[4c�P~Z�r�9�(R�([p��ަf[����gr���펚�ݮq�NJ�3��#g�Z���(s�s+�aKٜ�i}<"D�mG�`����^�4��g	�܀'��:UH�(�~�
g�� μ�s�g� �|ջqB���!�́�{ys���o �1A��+*���Z��#�e�k
��Fj�*�ەf��T�i�J�4-�f��/O%�����G��!uo�s��xՎƈ��o��ļ������Y]�Nf�@9y�؁~H؊�:��d��KZ�F���p��~��T|*��a�34��1���/��.��]k���� t!r�x��鑌"̮EN]ՆU���N� P�&皣_���N��
JlK�N��? ��J �}��$�U�Q��TZsV��I@��������[�q�/����|����+Z�lP����(�>8�>�{��&�U)�P��
-3W���h�����
qQ�d-�?0N"�5�o(�<���j�oe����2$��05�r����-;M�p+h荌A��w��Xn[��" �.�91/�V%��|�K�E�'ZFcY�>���E`��d���#�C��� �6+#���:~�D�>ܫ�kT���G�4.Y����I�����`�����߼K2\��e���-�̑]͒�=���~�t��h�2S4���#{�_,]&�����PB����H�߈�T8�uʣ�������W�AW���Vf^v ���ui�\���{����q�m��68
b�S�w7��� �:��D���?�{Ä����Og�Vݕ�-z�����9��J��PA�ͯ;M[�L���F3$Uքia[P>ʬ9H��)��=��ڍ$��`DT�1�m�͂��[��8	�3���vY\wQ�4<V�}5��-�;i�:�i M��U������g}�0�F�3�H|�_{&:}z�r����p��<�L�2{�
^ZC(V��Z���h����y��-��W�DJk�O���s����؞�L��Q���YF5�T��7j��}����ރ�\JPp��5�>����v�6#9���(l���20��Z�i�lr�����\ 9S�>9�{�C}S�o�7UrE�X��5~�:�\�ix@ퟐ��}�0D�z׀pWw�e[�qUurF�p)&k��IG�A�B}�]�^/Qr�k5;��aXMo��;ȊaG[��t3��Ӻ�6��ҵ"��_g�r���M:Y6f�HV����Uݴ{�֯E�dGVj3���+�Gn,�vL�TR��M4�k���0v���+Q��c�ۓ<gkPJ�z�0T��C�K��q5m���O#�R�pS"�*3����fh��ߕ8�s}��S�T��q).�rp�J`��x�꬀�wW`Y�ޣ6��������`d��&=]W��%�B7��/JM�ы�Rp9�\_1Ey�dC��ط��o�%*_S�r��=(�K��b,�VY�E�����!SϽ���a+u�Enᕍ}'G��CkE��rn���/(�J3[�����M__��&R�V
g��9C@�^�lL�xƓ%��N��O�齃>�#��>�h�䨕X��5�3v�/��yk�σY���e2'�S�2_�����`�(�\+0��1��1�CKO�G5�R��Ԏ�6���(!����79���\�a	=�Q|�4�h�x�~O����/�j+ q�##k,R9�����s`Pۇ�:�[V�7�H��O��^=���REF���n1�6��vY��GlQ�w��D}��Ϣ���,�w����0����[�۹��QP��9!x���#����������������W��%]� ��pa�|$ku/�������$�=ɗ'��K����N��T(_�G�Hq>^nd�a��H�^��{�b�Xq�E��q6�JTǳ8D,ԑQ�dQ5��)DѻdL��jm+���f��j:�g���/AܮP��X"pbĎ����5ަoJ�İV�~���u��9'P݇����RF�m��D�r{S�z٢��������9["5pD��b�W�WĨT�熦����4^eԨ�9�t�A/w ����+�%����1��B�9>6U�=X��7�R�_o�)�ڮ����&-��_����r�%ZU9�0���F�z�,�ɋ�<>2�?ϫYp��m�Bv�����< �l�[�1a˳�t�f?�[;�|���?�`7��]����.���H��&."d|��_8�nkJ��Dʤ"�G��,4A ��>}����[�~�6��{O2
a:g㝷���K�cU��r�s���.ʉ��R���BA(� ��̆Y��kI����{�s6҄x�1��Vf`j�(�Y-�����WN%�����o��A3�0s;}��ۙ��4R���D����̓���C���>Ħ���v%��*��M?�.��v�
4�1�{S�?gyE�����%�L�/�C��)��j�����v�Ρ���lv���_��uZ?Zζ�5}q�VY�iM^�&��J(½�T��+K�k?��	;T���IQ�~n��=Ď{�
ι�����#<��Q���RŹ�Oï7{uE������M�ưa"�ķ0��0�[°gA�(��1�oF;���to��a�&�>��Sm,N�47���xkg��f��