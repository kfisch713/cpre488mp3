XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��{�,�7����	 ul6�c벷gO5�Q�5��4絯 %�34�!k@��;��=��]_a�| �g@�c���Z�p"t)Oo�z���ݱ���d��'��7������"��U*[��><���p�/$Y2U��J}��[��5�+�C��x�_�0La9�u�cE�lÅ�w��P���Ov�i�B��>�IT��uS�4�k�5��Z�&e�D\���T?)mg( ��6ق,cNk���^^5O}�dcg������AΎ�3 Y�C�e���88=�#U�+g��9��'�/��Vhz�u�S��_zFDm�3aH �|AvUȘ�]�x������h���_�McX:���C!�j%��-��\�َ��֍�G}�C-��ע����>������2�x��	�%4�����U��?W��;��9�lg!�]�f�Æ]>UR�U!����xa]����N�P�"�rA�/�����I���I0y�U��z�X	[�Kg�Q~��i�M:%<b�����D�z�D�t��������;��|�q�$<���8��V�،p� %Fx�vG. =���j�4��e��R�Ea{�lue��G<������?�� ��&��Z�3*�C	Cy�H�H<��X�D�s
�F���X@5��➽WI��1�_x{�q�O��C��{fh,x��~��ۅ�h ���;i[J�*wv�C�$z{"%�7��Fɻj ��\Rq��w(@ee�>z�c� |���E�A(OK�:��H�k",�_HXlxVHYEB    1448     800DP�œ���7�����M�����ֿT���^�"�a��)��&�� H�?�Z��J@G�2K|��9�$�Uη��S~�0�ܯ�򽾶��e�����h�n�[���r��m�4��1���)�4LT,t�%�V�NhI�����l)+З���0�Ä:������	�%��L��U�44[����?�
Xf1;@|9�I}�&���`6x� �ߺ
1��E5k��ymx���L�1*�R�͇e4%�K��w7C��D�/-.��1��q�	X��o^��M�ث_ �8ف��ܾ�b�qӈB1$�0|#}I�w<
���]t��}�1a����3Fq-�wd�j�Cᅼ�I�m@x�X=���ZB��K+�t���,9I]>~9��Zɼ?}��ĝ�=r�	�ᦌJO7 �=u����?K_S��(��O�7�B"U�r�|�`�p��&���XhgW��&7Z4��6@\/%��c�$
�Yp��&a\�<ގV7�������4�L ����.�y���)�A�B��;��J@����T�Ws��r~���}��/7�F>ۂ��+��LMX�f�b|�b�R�N��KK&��W$Z�D�B�{rA_�9m���I�|2��d�b1~m��܍�{�J�Z���Sh��lQ)�kѧ�.�a���	����)}t4/[�
�i��E�H*�Z�ء���N��k���w6�K�o;QAF�ekYq_�;o8rW,TQ�b�-�5�LB��q#�b�l}a���#$%��=������C��1��gx�}ڴ|4�@a��bt��������!����6�-zS����uau�=���;.���F˺,��	Eޠ����P���Nժe��v�^�-!�B����b�E6�H,�v�p=��
����=�Cpϧ���6�k&k�3���	g���W�V%@F�[V�5�]��_��7K���Z�����'\Zf8��>z�.u�7� �-m��gm��A���V�Z��۲d<�
���}����hL��ʏEJ��u8�d�� cyI�v�;�YSv�;�6Nڃ;���׀�;�Zy�ާM�D�$:�/y�[�X���������pS+�Gi,V\'^���3��HT���D����e����0n���H����D�x��[E��L,���� ~�S���3ǒX��ݎ_w5���WOs~�c���t�P{g߈K��Y�;&�1�T�k����W,�"�i�B�0�ػ2Z�pn�q�3Q�wѹT�{��^��n����WD��7�3���~� ǬlQ��4\��y�_o�.�%�����??�o������F3�%��N/�q�W�u��}�H�KxVj�OGh�F���}KÁ[i�������֌	���򡇴utrO�CBb� �H�:�-<[��8�p?B?�����[�c��hM�Ec�mH����k�CN
Y�o���}S����y���'J��Μ3����۰/��'�O��f�④����E�E�Oöa�A&��F�EG�ЖP"�Y^u-�凭`�ò���"01�9g~�v��y��F�������ż|fwŧ�!�֟��*�y���(�猪�#3��]@)�e���JS
�'8�Tȵ��^ i��)b�i42��2�+�⯕K�V��CWﯴh�)*�9�P�
��I��61�~]�JGt�`,�g�\�^��p���Q.� %�XQ�|M6����l2G���X��m�����mW��cjO��tI/�q#5
�j�*�e%T��#y��4G��y@<�a|n\��M�Ʋ��#5eW�yF���*G�n��X�#���u!!v-s���������f�]����st�;J)���У�$ÿ6
��z~q��-��܇D��1͵PC�[32��.�B��J�M�y���C�}�x�!����v��[� ���$��;9/Az$���4���gk�廋��2lHǓ���MO�n_�CDQc�ꎱ`��Y�j��z9yЛ��	�,����O�F�ڧE�o�