XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��saj�*��>�Ð�������_��I[��Ix�uy^^�K%��B؎��pȳd��]�pH&y�"6q�]�C?��ڻ���z>��-� i���'�{^�ݫ&<��J��Q�rb$?��ߘt��_=��ә�2�9y�|����������g���
��v�+�YNں���@`ϴӾa�FH]˱��Ivhh0�1a�T�xv��u���g��P˿���i�h$*m�1�9
_������в��5pҿ̇��!�,�Y�U�p��(��yRqH�ڙQ�2-	��P��&0�u�>����~�+���C�QO"��$�?�� ��\�ot�.�9���*����_*�H �R-�����S��.M3̒���2�<���D�������v�����݀�����:'ڞն�zB��AH��O=Q~�|T�M��jѣ�ɒm0���U�_Y���£����]�/�kӌΔ!\�x�g���k0̞
���l������aCo#6ƹd�Ƥ����XdV�B���)����ZMx�YG���}c/�FYM0p2��$e���03�?-����g�d�oj�4z�l#���AVҩR�	���au�����9r�&��3n&n��컳�x��6=u��g.F(ZU�/�KS8+��>m�����.�Wq�e��,�6|��#�e'� ��#mm�&���9�P�٦sF�Ԧ�l`:ԤW��Vs
W[=�o�z���Nd=rQ���}�v�Ǥ�)F�#'5������bm �Z�L�gQ�����XlxVHYEB    4b9c    1300ӽ-޹�z��S�}�DMAS"���ߗ���"R�cE/S��F�NK�5�4`-K�#��<Ff+ul�;�&R �.��{5ʫDME�\�hBm-�/�>�U�²X��N�Zۂ�Q����e�,ϙա��N�8�/�h�uɻ�g�	�v����*)���m}m����cF��|?#��Ȱ	W�*��,��1�e>����
_��,�Zm�= �+� 搣���
�G��lu1��s�!��!���z���@L@��Z��o��n�EZFM<�=qe$���� �"�\$(t�_$va���o������)iq���Yy�Ep\UN��h�k���2�tj8�soZ��ˋ�#�����a�����w0>�-BP�P�AcY�9�8����+��;�j�F�5��3�on���B6���i�d�6a�tvs)��5�I���HN�Y�H�G�Y��k�!9��j)���[�Mu�~e��k�e�F��`����Ұ|!�����L�8�� ��].�2�0�Yd��ˇ�6���D��tU��"�5��
|�Ւa����t"-�/�:,�>�L�a���!��S����$k���6>~���=��֩0(Oג1�+��1Dc�a��dO��/j�ݚj���;�i�����@8�Bd$��Y���uF���r��6������#v��W=�-�l��+/gsV=�<M5n��
��y}TuU���t8q1'L��Cek�I(����1����W��#m�ήk����9���snXv�KB��!�[:aL������
^*���Ei���D�R���ޭ��F���t�<$I8n�{���:Ѥ��O2�6P7<{��04��rQ0�v��~�������92��ۜ���������9���+��z��7�d{H�x��\�`GH��5gȕ���IcE�Z�b��/��NМ37,��T=�*��[GH�����´�])t��i�j(�;i�!!�2%4Y	$�Jg�; 4-萋?��r%�<0�m��E����r�/}֭0Z O��������t¸�mo��1|W�Ǐ�1nj	�1�����bj���a��-��N������s�o�dc,�r)�܁��H����vfH�`2��|"�Csz��_@��(le�a���R�O�B�s���'8ĆjL\8�J
��]���Z�vu|4'�z N`����P6�����&W�����N�y�t�������!KӬ5��Z��m�����s1/�A����������v�������_*
�jd,�Q_���߆��ʮ���'��&�"�y�s�K����G]���+�\nk�Ihp�:c�e�!$�"�)w���9d�����>�:\ls�o}���}��Boā�N��K��#�X��p��q�|�X�@�F��u��1	�X��:���S�3?����i77]�%�"����׳ZL�DY�3� a>MZ<��(��y�)=q#�U���1�f�c��\r1Ջ�����h&+��u���.�#6n��z5��{��C���Uq#1q�m܃Ҡ�������N9�����1G�2���NȾ����Ҫ����j,Z@ d�b��,"�z�*D�\B*i<pD�ۚ��c#ﺌ��ڞ�8�< ���%�=OWCl�`2��f�K�+��$7Y|���{�1��p����det�=�Ɇ?�ٿ���oA���gt���Z{:�d$	��Y���K��X�S�� �2h1�M3F��BL��XVϜq}cR�f�?��P_��/*W�����R �`��Л�[ɋt2� �p_%��}�k�����tV:���E�
=P��)T�~>*�a��*��>ѝD �z�q w�VN�D+O���#�B��B�l�-�u��(���&��T���B�Z������CKv�Q���G�2�V���ӏZ!-bTW��;�������j�b:k��ww�yKs:�5V�+ؓ��l�OK]BSW&|6�[�,.�D��æ����K�0F��jT)��^��J7$u7-�۲�:~�I���?��S�P��a�u_���q>����3��.4H5J$�\Vo�;Z���M�=u�x�U{�"�9h�N��v�;�s?]�U�v�b�[�5�[����ہ����aD��o�T �+.� ?���Im7q�{��i3���(k'� ꎓ��[8���r������?���h�! w2�DO<�cpe:*͢��3� M	)� �$��p�#NyjD�%	E'�I�Rߑ�޸��"|z"O�����t�dp@�"��jr%��@٫>�閔Xx+-7�����W˾e����#ڈ�rn����K�L,Cf����6���TE׷���#�;��}�S` ߍ���Ex������R�[�P;p�i)�����m$ ��a�L,ixo)=�1�W:]�ۊ��#������8uYZ2�IF9�]��J9#͈@���yx A���~�"Ev`�xT�-�PY �JVB�ЇIXC���`S�+|o��Ǝw ��m�����^Y�����is�M�+i+��TTV���W�-��7��KX�^��
��m鞁Cl�gרU��F��зG�*U�w�jgл�r�6
hcG�����J�ZV�l��V�����
y6r��Z�\�J$.f9��I=qC�X�H�v��j�W1���;�`�]�&����^���x�mF���˕ڀ�;2�i��|%h{��C���ّq�i$[�N#Y����<W�G�5$͉�;թģG�/N+�]�P���]���u��Z|o�G~3�$���x�q)sK80�<�v�Mfi���H��w��8ȡ"Pq�α.V^[��m�v&�6{���rX����qK�\R��UI	ȡ)�Λ�6�ܪ�j��>��=R���w�w~_�9�ҋ�`��3v�KJ�Z��HӇ���!����*wX+�.Ȯrun��h�R��>N�Y�%�)�o_��GHuL�昄�oD��HmG�MW� ?�D(��e���Ur�S�J����w˛�Ȕ7y�4XPN�䰰$�7L#B8AZp�n[n��i?�T{5e��%�_q����Qz���3��4�F��_�p���B��״ߤ�գ��e�fk�
������+�G�"�L��Y��L]��=�@�����`5~�P���8��#&E<\�FK�CE�v��bX@���� c�V�����w�`fJ�`����(����v���P�PFv�1 �LK1����#c�yj�%�&�T���7����l��"�:���r�������ѕ�9Bx&: q�Z���6�V��]9���ƕ��U��3/�J����&4W�(�pP=@_��tɠT��+ZY����֑�g5l��g��'Sf�;Q�Zpc�W��,<���+
�K������Dɤ�0	�B%�X{�`ȢVb��C�o�[�h�&�|`������;����'� �m���yw;���d<W6־H�����,���6� u[�<b���k�zg���d��<gtaA����b�W/$S�>*�-�[N�֚IR�jp������&1�H_��
�2w2w~�����A���=M��!��g��
�Ö�.<��%EӁ/'������|:,��r;���ƃ4EJ�b�O��e*H@0����[��z�>ӛT��8V����P�����⁮e~���?ؼ�b	}�o�N���%J>�?��ӂ�~,�o�h:��N����{n5#^���ȭ>êC�*f8�l�I�l;�v3)u��l��Df��!�
_�F5ꮿY�z�-����*h��<�u�2T�]�K�7R@X4�{x��ɔ:�1^���e�����m�:&�Ք
\��a���>� ����|%3�T�7��P����h� <Bx�tTB�TmCtҬb��O�/�.=^�e����Q�ޖL���U�GX@�	�kMԌb��V�<��MZ��l#��z���0��Ab�@�h���u+9��h��`����93l��������B-
�?(�g��?�#��^@�F�GUڼ������H'5�"SW��m�r<��:�3x=zG�U9���~�l.{��9N�B�a�k�<x�rF����i�W����� л>M��/*8+$s0���i��Z��^v]V�\��l���<��^��;V���A|E�Ś ��1u�:��aEM4�K9�5����U��;�)�-�v������<noqY�v9��LO��O2h���9N��}�~+eB��Osr�6��j7
�׌�&�д��?�����X������a ��4`O-�0d8KC�|n=�.�������؋���5���8���L͈u��pX��`A��ݸ��r0�b�3.�~oT����!&�����O���߷�C�v|�S?�J�i��qs$���Ih:�ۗa�ޞ>��L|��Boh5�ڄ3>yu����ˠ��-\�l�<
D�:�<8[��::����>~p�MK]�n:+���%�'K����~;��h�M��~˝� *�΍��� ��/��{ES�4�)�@LOsBlQ/d[��l4�q��)+	�u�b��Wh�O�/�'���˺�ݜLӾ���pa-�G������F
�fN{����VL@�%�fz��i>��y�A��]��p{�۠Y����pL���d�
{��x��.ݯ2帜^����`���"GNVnB��)�lf�
ᅝ�s3Qa���3<�)�G�D-�B� ������]�ٳY �g��3n�v{��n8!����