XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���i�(ڎ䍱����I�B�X��˲�IMt���j��/H$�<����_������#R��P�
�ĭ��+)�/ʰB�/~c���\R�[K�n�;��KTe;:T	�N�NUsM�?�wt��Ԣ��j&�Nw|Ct-�g�dT�B�z�8f³1�����$��T �i"w� s�`���uC����Z�pв&'� $�"/�&c�4<P�=�q�<W��0Gg[L)�O����Z�(�6�8]����I	�R�b�����jk�#�3{�h�##�#��'舦�͋�P4#b�S"E�U�~�j��ܾN !D؎8�%~��Af��[�JI�k�Y0N=����k�tI��{���]aC��6m�D�.��6N�Aߺ�J����	� �Q���t��WpFCE�$�@dU^���~���A*�P܌e -#�J_�Hs�$k4(r��U���%�(x���R��u�#bض�s�3rq!u������2�H7v�~�*x�g�@�?r��璘��ʍ�O��^�1��(����A���ߕ�6��� AI�dV�	�<>���Q�O�R'�	�F �Қ�L,el��6%�e�5|��3+����;,��®z�ʼ:ՙ�z����
&�Dr�m������X�mn�1�|����m�B�Z�������P���~uA9��s��q�� δ4����~�%�>�u�[���ɩ��H5
 �P�#6zS��se.}Ѐ�%�kX�{�A�.�ܖz,�Z�f}/kXlxVHYEB    241a     ad0���C��̪$���Qh� rwf���1ʈ8V�)F��[$�驯�zZ�f�UDdx��͙X/L�4<ǀX�F"�@1�����ƕ�Ṕ3O�$iU�\f��&.�lۥ��v�����>+�ϺF��j����]���qR���f�uβooe���c�oWnc�K	�i����r50�q���C���5����
����/�X��Q���Ӝ.t��k�1v��� A[�����3u�gw�j��W$o�j����S�]x	{��vL�*��_Â�B잎���!�c�%T���c��*����?�N�xy�7�)j�д���{ �^����G[P);���g͈|��1V���	��ГWnp�at�������Gohp���f�L��� �^y�o�g\ ;� n�Ƌ9�₼��m���1B�����ށ%<��^WT��X���Ǆљ��q�dg�-���sB�uDV��n]��Q��ۗ�b>x�^"��͸�om&��p��b61��e�M�asK���Y���M\����f<�cW�/2��N�� j7|M��'���h@����P����(��qZE�ڂ(y����H��(�gL��l<�� �i5ۍ����N2�Q&�jP櫧-�d��5(�7�Rx@Y��n�Ƭp�=��}�p\��b7�n�?���d�'OqxT����\«� ąI�pM{ħؔ�o8
��͵��*�4�:{��vT�5>Ձ#u�{�����9QB���ͭ(��b]c�Q�kb#A=HJ˥�?�pw<�� �!2�7���W�-�����{Z3�y�)jq⣜�ɓF6}8_����	8V
PN�Ia��#���dHDX��.�RRW��y�}qag�U�y� N9�'\����7�zl��}�z��W5xb9
i���r���̾6	���01�ng�ԝ�O﹖��ȍ��֟�9")u;�eF}��ar�</����E{'���B�[���q�k]�'���{F�%n�L���P}���r'O^�
�$4�&�D�cN��Jף��&9CF��� �$��No�A���V���DG9v��v>Tvα�}<<��?ݏ@r��]�!�Q	kܗY��G?_�g\NZ��'sϕ���{����g���&vw�*�y�\����2(�]�iy!�s ��2��ڋ��A���BǛ{��,o�3� E=q�$��v���dMn�7~ɝ(g�(4Q��[c�d�:�����IN���%�az�>8�2��w�[�wr��1�dg*�����*�������[��ߗ*ic�$`'ZA�݇=&�3���t�� ��f��K���_�>��_����-�2���*���C�����H�r4RC[G���#�Z����!@k��JlJ6L(E ��(����}�k�g�7�W�Z0�P{�P���t��M�����B@�hin^�: ���7��1�X��k+�X��c"�)���b9h�p��"��F֢(e�&��^Jv6=;� ͩ�Nq��������Jz\3�C����<��h"�y������x�3����㙴�kQs�rFx{�^��*C��P�Q[��*�v����Da��8:_�5�,���R�	�h��V�y:�M�i٦o�nt����W�9{݂D�y�@js>W�1>���_��{Ou��7��إ�N[�"F6���J����E��w,��vv��<��oe�y�¦�9�r��;�!����/D���?���}��k�Y�X��`"�@����'���M}�5���j=�;��T���	]��ɂ����o��I]M@���v��ϑZ�%|�(��j��A�RC�LXG����9�ڨ8�M6y����M�0�F�-迍0��Lxp=�6�@(hխ�`{`�.��X(�g��A_���gX���B�5-|���Y��y#d�m���[{�"�6��+$��o�Q����r���:]
��.����a�)	��ا�����w���d��0З2�fX��3ꈢ{q�M���u��q��5ڄ^ {��q���%��Nh"�g������h˞X~�Iϴ��\}[Eˇ�ۯ��}��4��3�TSa�D&$峽��.��0U�xg��ԃ���Ola��Qa��FV�#���0��� q1x�8zw�ml��u&^��`��e/��g
��Q�n4x���iЛ��Y&���M2��I'�����; 0�\��MdM'f�f�c�������hU� �&+%�şn�dU�״��P����y������� �maU��d5e\l�Is0��r��1w��X�cc1^��|C�M"C��ɽx��m6�p%ꬤ�ŤX��mg�Y��Y�a��ݣ��@��WBzJ��,V�E{���[�J����?М_,z[����1��f�J?��J|���������nn�g���5�pI���F�wo!.�Cp�kֱ��K�s(=�R�Q�f5�p*��vI� �!ooܬrj�`��i�|��)~,ީ5vgKk���8]�ě��'���`��3��ţ����8�Op�����?���u��Խ��U���(�{�"K!"D��e�$�b�ߢۢ"��P-�*�}���%�}��r���`�x�M\$��b�Tu�0t-. ?��S��M���%:���B���O�@9�̿C��|�\vX�g8��	kAP6�ƅ�2����������f���/U�H:��k9�N�'����D��~nG��El��W�@��VT�