XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��d��\�C��V(��k��Afv$Q�����3L�ƨ���# �a��ip~j��u1���f���Q�7{��$�'	x];پDU���9GI���^m�x������em��ɡ֭��ɻ�A�b7�~���Tߓ$��	Ĩ�)o��'6����1&y��`�����WH��5���Vq�7>+x^a�5:uI[���p�M��#�z���*���2��(�Iٳqi�&Gbs��M��r�2j�d��X���>�q��\��?�~po�E�&u;����ؙ�>�d%':�@{\�c�_e�֕[*IvP�Y�|_��{v���>c�V�.E�V�y} `8=;�����t�O�S�b?ޔ���f�E���W3�Y'�{��?�9���T��<JC�#���K�2�������%֫]��G��ȱ	hф���F=ug�*�����4�( �?B�Yu[�*2U?���~�O0E<N�* ��&�V������ߨ�Ԗf�"�bJ&��o��B.�gb�z�X�Y��$�!Ǳw�ȤI*��uS�~��gZθ:̾ڴ����ر!/��χ;FX�*O�E{=�-$l!#�k���<�m�D� �-�}4q�.�� 8����#��jC>=��:mB���&@�R����=G3*@���ipt�0js�V�δe}����ţ�^�n�Q�f?X4�;&�8������F&� x��P68*�U�;�ߋ��"��[�-�����T+kU0��j�m��+j��.{~�ʪ���*XlxVHYEB    1a34     990�"��^c����c�Y>�)����?��+�#����H]�?r�hG��np�԰:�!��5+���t`��1K�f}��1��5��ZhAv��c��l����^A��G��%Q������@�K�3�����g�N�!���]��n��fo�	��?D�=U�1��}�D��q�R�c�K��}&}"?G8�ܴ�h���g���D�6�y��1��&mYs�6�ȠSV��-�[(Ԍ�D�g���)� uݱK�o�L��#H,�yykJ���4�L��2�R��"���I��,"�p�ըXՇ�y��~��@;[�-��� ��K8����M�=�Ƴ�L(���!6����� 85�JfM~qk)��5��<0Uk �uǓ*�{�k������3�M�?i�I����iaɆ<�\�9�	�A���7{3/Z�}��g�d$y�/�׿2����z�:z��F���rn}��jz���˔(Y�1.�+���
��Ŕ�S%/~�Cw/k�H?
�K�R6)C�E��r�V��P��cy?Ŗb-�k��7����#o��g-�sF�<�h�Pg2X�3��rR�:m&ˊy�V9�g������BeEڬ:Wra��_�h��P�V_žrY*ݲ�<)b����:�#)
��"�[&ool��F��1}�.3��:�=|c�i�qCU�}B�{B��#��ma�2��sk5�6*��� ���eK�/vd o�����5P$߀��0���2�eq��;@����ҧ�Ha	�zh�%��y2����
ө!y����d�1�#�f�Q��a'�_�I����}���=�6�ܺ�xL�����ѐSOD۸�@�/l���?�ݘ��XŊ�7{��G��Ȓy~ݢ���FcN�	zY�.�,��g
�Cݺ����_e�,^Fi�{}�c�t��6B#�i��S����b��b��=�U��e�Ǿ̠��AIw��p��Ed�dkY��w��Z�;bvM�c�Z�Ⱥ~�#C	%�J�y�H����#��zPd��})��ф'��&��m�ZwQu�&�2��6���Һ�;����ƫ�t㌫'�R�ɳ�ͅ���T<q��J3Y�ڸ0ַJ�D(�����,����V._%��R]*r��8L�m������::-y��(�\Z��I'�aH�2bB����9߲?�X�����1��W���BLo�)�:]�'`�;���l2�M�I)ؗ	� )��;:��l?��P���T\P�� zt��Z�Sa:e���}s]_R�dM�#"p�N���
[�Z\n�߭�|�N�L2HS�*���};�Ȗ���Z��V�� W�	H>@����� ����2	%2Z!��q��G� z>�'��÷7���U	�(���yfc�[-�U�O~P�W9VF�����@�ry�(��`�/��=�����yG��}Q�~��M���~�=9����ͽSŬ:3M�x>\��jnMg���56!��.���k�9�9�n�]A����Ց�F����Q�ܨ�B�<��2�W)W7�[J�5�Б���`c��1��W�4`�$�ԙʃx��F4�5�p;3�����WbK�S��7��l�C]���<�N��0��f�Z��Nj��B��8eŽ:_�U�v�ߠ���r_\:��+K�A"�d$�Gf^��uL�V�>��?yk?k�7�1��|�����G�q�b�2���g�b���ׁ3 ��DbQ�W�d�l�����ߞK�Y����f����C�zC
�pUs��F	Y�L!vx��VG�mq�P�k�ټ3�VTJ埫�Gg����(U��lu��0�x)2Es�������w@�3��[�~�b�ǅR�v2�uU��x��0���E~��w�,���~5��DƁJ��/��"}!li�һj�5�	B�Q�s�O�R��D�<�{��p��)��4�~���՝�Vy%���§��ȻV^ų� ����Ē��h��?��t�
��X�)G��IXoE"{����: �Od	r���`��`v9�[� L4|,q���Jº��Bl,3�/y��Fb�
���.Rj:pw���yâލ��n>�.���Ñ�������t�]�º?����/�6�܋��<��5�0��v�g4�J0�!t�ҳ������崣�4�>���LD�����F+-g`�-���F������ l'W{)>���[�LDd=�6��u��?��S(�"���_���36 ѕ�b�M�8>*��]9��j������r{!�"Ɇ���(�Fw9fǡ��Z4���ʥ��<��t:I�h�,]������-6k��;���/�=��1?�uf����W\��%~�n�j����!2D��{*Vx��P�U�Y	�7��5���Po�	h�pbk�Q�9��˔���u�&�/h��N�f����}~٨z���O�z�5oST