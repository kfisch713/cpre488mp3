XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���vH��ߔ4��1mO$���kԄJ����5گڑ_�
X��RΆ2t��w��f�]�9�w�<1^�g��˯�9�L�o#��4���~�s�ͻ"���}nm��a���r��YL'=r��i�]�{�����T.y�xY"U�|B�*��*�J�d��R\R�F?b�[%:F�͝�ۆ�ӫ^p����(�c�{��MĪF<%��_���=��������{��.�0wc���[D�4kz����;̢g�?�'x36�ss�e��Ak#slc�*M����������$�^��(@�>ԽN#g�ec�f��<xH�R1�L]~x�(�HK�@/f�E��P�k�H� G�5�V!v��{�t������@գ�c{ʍ�b^�dЫ����MWó�����+�� ��f����dt��UJewH�˴�0c6���h�)�5��.�\�?d�=f��lY����l4���G�I�'���J*6�"��g��`��,�ܵ�PB����	 h=���-)�u�wN��ȯ�4Rtdm��35doD< $c��4\Q���;���C���^@�K�&sA��Z�g��7nQ�{�P�Xvp����i�<M��2�����c�!����e�[䂙����D�X_kt�-�R��r�j��(*#l�5S3ܟm�1w�;�9{���4Z��y{'17�Ϟr��LL�όw̺=A��������vI�.�M%� N��A�U.�(�X~�2v`5\{�b�8����:�S��XlxVHYEB    48e3     e00
�k��zXWPS��J�U�lf;_�*��z)V�:1w��PM�B�N����U��݆e�Jۺ�-KO�c��k�8KW�s�2+��ѧCB���$�C�#�u�և�)�[�X��%�$@��e�ы��j�m7�D�7��+A8����R�h�]�5�hA1u	Sd�S�r r�f��=�PռM�[��d|8u��z��V�B�X���?_M��TC��f��PMw��`L��,�XfL�V���y��^�K�Lv��V�?�r�F�F�
�����T(�ve#cD)����]Ab���R�$c���u����"���RZ6F��E�L؅N�cD�{H���sw�hmM��b�Ԛ_�O�����R�y��h�m��<�F��B�㦥\A�>z5�ᡎ�L?�U�7(�L+_[���r�;�������[�{=�M;��=��c�Zg.��Q݇h���xdf����}~�8�Q0����w�+ʸ�N��S�Բ�k1�oą:�1/�W
K��}H�oy!�]!k���Ό�n��Z�l��|�#�j���g�z���JeM��'W���6M
.Fɂ�:�׷o<�<m��ߠs�ꟷxH��V|x�6`�t㤞�����M{�T���8� wO-4!W`��,��OW<�QFr�x�pe�X��6оȾ�ڴN�.>��{�z�� ϡit<&Z�����	��l*��C�ؒ�w򶅯������b�ǈ�ᡄ]lZ]	���
Z�)� mڑ2���1�5x
aok���:�Q�|�J�լ�dn5�6¯��(h*��}8o��"��.��j�}���véՏYJ��b��:�oƻ��aZ�~�z�Q����u-.�)�O�k!��8S�A@˗T� U���G�~ޱKw/�4ډ���͏�n���gX�/Yn����|k&#��MW�R�\���Lv��}�>SG�}���.���wY4�׃�]��3�ʃ����#��!��9B	
2���J�<�Yqp۬�n�Z��̖I���BG�8�Y��.]g^��	�v�����0�.y���Z� �p�=,��+^�����v0`d]Y-2����}ʪMͿ`�a;m��b�j���@�#�[r	LU���]H��.*��e��f�+t(Ñ�˿���\�����������3�nDIa�,6��$�h n)��S�h���oK�.����������,��P��2)��a��h�{�
��T<��3u^�'�Xlnt��
-7�	�ӊ�62��:��"�f�\�Q���h&�.KM7�����l�|�}� j,e@�鿰�Y�/�`�Fԣ?K����\�"�ը�5
g)<������k��I����^z ��y��?l@5���C���*,�8nO_��!^�[��O:7��"��b���N5c(��pW��T��w�^[���I����2���O��ꦧ��ss�d��$�_��u㲯���B��Y�O:j+�}�6T�<<Q`�3�w��؊�e���!VzE�ߵ����wv��E|�VVp���3�B��|� Zv�Э����O����mz�Y�58��`\�)��}����i�+�= ��n�b��C���b�������9D ����p���{%VX��z�ef�� ���"[GyM���dȎUkL�@�֡W)"DL�VuCouK���œp�I�⦂��M�x�j�Q���oa�HҶ�~�)��R�\h�0�p����e����+u 8[�<ƛ��bS
�g~y�5��1Ҭ��S��^�n����t,�c��yu��`���-v��)�'���Y�cl;a[�5_GO�с�_�J) ����c�j�G����0�^ґZ��b� [S�;=[�0�ʩ`�@7rq�fj��/6^�-�!��qk��"�XPB�%�?�nL {l\�ykѾ��\۪p8�̶��A�l%Y�!����GBNځ��ZoS�_g��R��'b�)#D��$�Q�� �*^���8�J��͊B9��!:�JI���� l9�0�yB��d�l���Nݯ���o�1��>�0�{JS�*���t�oM��C�� %
�O��%�Q]E}C��B��C��$W����S���K�<�	X����]��.��U��|�7e��!�-戄x͖�/�Ʃ^�y�s��~������/;��o�jշ-�Ȓ)���I�5���e���\�������u�'��|�X�t��	����՜��Jh�D�U�P��K���롂'p��Ι�cvo�����J6����Z������1X8<���kuwW3�⥙����o��������&���u�W|�5�;�hסB�ֈӮ��^��r��^/j�W����RH��~�,��*����mi��� N?�5fP>^�%��eo�{;���br�"nuh�,�ɮ�T`�-�sX���8z�Kw�uphɦV)30%w�Is><@A���cl�R���e"F���|f�g�����Ʌt�O;=V��NN܋�w�~�hlH���5I�}� 8���n)�Wj)�����n.�P^�z�FC<k�0-��~���!L\�>-8��}���?x������:���+Г"H7J�Q�����i�m�W�	/���y�����j��!o��#W)x۫1��'��?�X?�Q�fxQ� Zϓ#�B�3�pO���t��i��WV��
9�^�˺��1O�)^��4E�����A�'���vK*3��}�+�G7�d�Ԧ�;�!�F�- ã�`�ӛOC�� �)�ҝ�B�'J�_�ɦ�y��l�˭���l!qN�˸��̍+kA��P 9�X�fu��.ٌ��3��f]��R�2&,��aL&�4 q�TD^�����4�s{���H�#�)����(�2t4G�I�M3FT8[d�L�A(�B��>#S/�W8I�T��`D���Is�L,�Ô!�� ߡd���!��L���o�,A�t{�X���x�@#�����?z�of�[e��C@<��=��e���Y����Yl�27�Р�4��}5Ӯ
���:�.��\�O]����]Q>hǛ_���iZ��)���f���`���6�#z�������¼����r�Y�V��ӯ��o,�y	��~k6�$��hHԘ�����Ϣ�5DKA�#��<�-1G\t(��eT�5�v�z{ko���7.c�{MbS�=�=2�O8�#NТ��B['D���Y��O�� ��otR���#�t#�%,�'��}ȬFTr!��tXH�	�S����~SA���@ ��|$��86}��:c����Yt���[*Z�WjL�]<�⨉󾫯��.��#���̏=g5�>^��Hحի������-�6�K���S�;�U�%�;8r���^LA�6���Ǫ�����k8�ɂ��<ʓ���6�h�@Ñ���W���m��V�I�=�,���]��}�(��o3���]�?M�pS?�i&L�|V<��������WF9���>�!bS+ ����T`!�,{��