XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����|q��U~���c=��ț���A�a���b2r��c��d�����z���rL�3Er]/T^�����p�_��}V?��C�����zκy��+��1��5jP�Ͽ3����&��/h�^A܆a�v��uz�0�*(=V�VZ���孓�^��i�R
�\
Ր��4c�v������i����4���FA�6�º��+|=ݬ�j-�w/%��ZHd2m״<�o�kd�D�9)z�Dμ��ǆ����җH��aoh|1��|�-6��Y���Ϊh��h����L��$2I{9Z5=):M���y� �ͧ!�t�l9a��:)��p�����4�MG��2�2S��gٕ1�8ݍג�]�%_fG~� �*�W,Τ��E՛�V��"�b�H?�����E�Nl�,#�`�T<�%�x�{%�������ލ�Ɲ�4j�6�U.J��o�^x�=罛-��R��9������n�Xl�1m7���'*K�F14<�-�6�VZ(��Z��m�|�,f�`)��7��eÃ:�q2�b2�g�aq]49	VL����w겆�А�I� I�{( i]�S@B��0�ŘN��E�ed�(�wm1����`\RU~Nx��:߹�;����$��3	���~���A�������бO�����,����Ɂ���7�U�;g�� �Cq�/���,j���U+ C(|$h�ؕ�r�7���ҧ���DO��'���e��k�]ʄJ-�Uq�āgi����61��7��C�}���-���XlxVHYEB    9fc7    1fd0�L����Xs�̐�UM�Y�ڡ�s\y1
_㊶�������r&|<1Z#>*�<���E������^�P�L+0�f�����tD��4�(�!8�Ov�r��,�*�ȵ�%�����`'vW�u���4����Ӊ�%=�A�YCۦ�p�����E��ysWX��Y%GPp�c!�taZA+�I�N����ٲ~���vR������ݥ	�!�DZ�8���_�vb��;֕�K^N���n�1��ӥ�L�ޓ2H��I��ns�HB�K=C��W�a�����Vo������CQV�-�V�(�R�B,�q�o���}��)�W��W�E���/7��B`�8�J��ʕL��n��Q��N��M��w�I�%՗���V/0h��@����ݷ�b����%�iJ�B��8h���J��ȍv�r��\�P�ǹXa��i�l�W��.ڭj�RZ��98�kd�q��~ַaeˋi��0���D�IK��"u��'jW���c���YuNm�j2@z����^��Y}��b̺�Z��+-c�v#G�a��Dy�������]���Q$���`��4���B����z��J���D:���]�N� .�&j
�4 fdU.���������AH���m`gF"B��;^�9���2A�����z |��W��[B����&�����TI�z�l�6��C�����́FPp�� kv?�7�2�Q`/���^���A_HPO��ݸ_>[�#�_@╱�Q������v^elU�J~�fᕚ2����P�2k�,�̎�u��W4o7jdo;L���'Kw�"\$*V�����,�]�T��r7eI�"�2�yy�N���X�ǲ�a���y�{�Z@�y�ɏ���Σw��	�&�Ո�IQ��b2��'T�< �@ i�S`��=D�n*��5�.ǶW�ܳ����dd!vd ����"�ҋL�{?�I>�@:�I�n��H�)?���N� n��F��yg��`�.^H��;}�H���o�=���;���I�yEW����y\¶�e��y�	1�X���t۹���\��`T�w�n��#��pn`�6b�o���:LI|�C�Q����n�gƛX��?��]��䱺Ўi&>969x����=�7V��q6}Y�~r�=�ea�y���j��9x'g��hc�]Ԡ���Ѓ�����=���f�PI��pw�
�p�`^��NL����񊸖�e�,�?V�Ҝ0_=���F��j:�xb��뎹�w���2�0��{�EMR�ͩ��&��uG���u��b�����퍾P�RL*�+�i��oOy����2k2dt�Ô�vp�k)W��Y�h�����r�Y�z�O(�i=��N�Y4�y������w�g�:ll�2^�P�
���3��A%�Az���])L�ZT��^ݻ�\����ҧePl��*#%���3c{v�U�)����Ҽ*D`u����N��{a\X�L�NT����t�,M�uo�_�\`IU�V�}$T[s,ٰ�M#5<��?�d��L�9է6Sa�%>a�8F��LZW�I����{Lw�X����,��i��cn��5xP~�=�V����Lx��X��-0C�����;������Ѱ?i��q�
;�d'O�����8a/�(r��R��5Aq���7 A���*ڸ	_���U��c�U˿�c4�S�l �,�KJ�݄�:rg��E9]�U#�b��w�ѷD~��.�H�7}��Vb"�p�gő8��D�ٶ���u&
��A���%��ղ}-�Q���vʱ��h���gc����R�΁;���ꬰ�_yC�W�Ce�!L�����+����-D�ŵ��E��'^�1]�6&з�f�c�t�,���q��������;#� ہǟd�<���t�O�������Ŝ\�U�;�uܸ��#�f�����!B�ٳқ]���hE���@�{-��v�+��|�2pj�EA��6r5WAQ��Z,�*��3���x"<�JՔI�Sv�����*��5�gr�+�È���`8pV�F�*=FR�G�O KX���0]Ą�@�/t�5�[��'Q��.����|w���~�n{�$w��g#��'b��A���d!���x���:<�.�f`iB���(����1��E�<���rט�M;}(��S�����i�J��<��$���<x�����ڸf͓1��J�k��A��XF�C�
�9ߛ�0M4h1������6��L����K�.�p�Z�Y�͝�����y��������q��5��!w�m9�w*��n���[/f��<~�����0y��~}�ER?��3��ke74�Y~�vi-�R�{C��r�^����%�R`�&Q�qR_����� � ������v����(�/-}�a�q¡'o*q�İ0�Yb���M/3w��e�b�L����&N�*4&�7�!�g�$��>:�dh�TW�
�&9l\�����kc�<qmJ���b�*�T��$��ݭ�y��|Cø�7&��2��?,(Lh�� g�=���M�^%,��S3>x�mZV���הڽ�ǆ����VO������ɬ� cߜ:@[4'/�i�E��e��7�o�#Y�H߫�(��Ү�KOY�	8��
	�*��g��Х�#C�7�ԃ�0��H`��%-ؚ���A�+�;s���498�Иe{O�O�]u�}U�X2+s��Y�SJ��9Ƕo�&��S��^�Z���֞�ŵ�n�����wMM�Z�/�� lݽ1Ib��/sGxV�(�}���л]2���TЁ1�ss�εQָ8GCUc�]�ycG�w����'ar��y!�Zlt�"��Sn��I�#�U<��k;R�='��Vzq$R����=������CLf���$Tm�1U�Xi8Hge�]�M���%�Ӂ �
�y׫��1c!mb����lW,�+��"�I�c~C�jM��vx����x��9fHM?�w�ۆl�#3��d��a�мi�����iG9���C���j5n�����1�#���wy��P���^��d�h��W�A��'q�{x֦D0OѶ����#gon{�[^\9��h������㎞x�Kf��V����p
�F�9�:q���-v������'���$C������
� �R�I[��/Z640!Tr��5���8M�������{Ug7�뭼�|�^e{�&�Ax'�ݫ���g����� ��A58;W@��g�/A��r>�6�}�VA�D^���21ښ�0DZx�
��c]��c��9��̴���,v�Fs����
ZXPs��+e�qSJ�l�xԦ����$� eCQ[t[>�-1��SSi�V27�D�������G��ˢK#'������&��N�XuB�Z$����jq[%KP�d�
{vVh#$����6�� �N^*��q����ҋ���X�R�˗�h�g2P?��D�"n�݁r{(�p�l�c��p2�Ș�"�J]�:����J���	ȳW��)�����h7(T_ŧ7)j����nwhc���))q�a�!���ы���	TEF~��]��a��AFH�p�0�P�+�H=A~x��fItq.�v��0���'����p�P��3�*q:W���,�������P
� j:1yp�2��u���KW�Y�	h=._��ڼK�-�`�ޅZ�cck���A�b	�Yn���{�����>�,��S�#� ��V��MГ�*�nf���r�	H���D]�X�9E&-�D����c�v4��W\B�4SB�J���.2��S�H^�P����$%���T�^EP,��.,`���a��o��f\�x�W��o�" y'y.���v���۲31L��,��"˴�b���V�-��e�ZM˞ps��gk�{���ϭ�BAJ��$�C&�`�'��%7��f}o%샲�5�j���qw����'�������w�� �z b�Cp�I�HmY�X�-�1�v���G׮5uD��@���iѺ.����aPc�߸��9�l�����0?=�zR��x�o=�ۨ*�,�P�b}X�
%���n

7FNZ.�1�ʒu�,��$)}X�t3���s��0���ۻ��|����\f��y�;V�h�����>�6��Ժ4*K�l�<�xf�iQ�BP��@��\?ڳ���;BϺ'�ر�L٫?LJ>)Rw2<#����3���\������|帊o�ahf��l�F�P�YZv�	K�|_�z�L����V�0���p�BA����x�;X�:L
���mOϳ�/q��0?�l]x�+(�Q1�L#����I�AЬƎ�RfJKd�+zu���7���7{�5�ⵆ��¶�B8Qbi�Q����hì4G]du�%,$���x�L��܀Q����G8$h�(�T��H�I�F��n ϓ���3���|�q��R}�!�; FM�L��c����KT���׽����`�:#�w�	�hI��-j��M�)�����\�4R��@.5w��LC���AX?2��v���.�E�L�w�^�����S�(^׮��"��K��(��~0�"�o�f_]^�M��P5R�,hM�uԧ�����b���f��]l۸*lFgUk��ň=�������P��i�+��C|Y��v�۾�A5�]���"6L��f�:}>d{����=�&�&AX�Q�������Q?�QH��ZL��A3�	�� �GTA�<	/�ɢIx��O�a�?�Bw"��@�9w�b@pCdxW�vSȃ��[p��ye�w>z5;�T�Bp�P�N��dypעa VI������������7 =���J���;�yK�Ѹ���v3b��g���&������y��lA���� �H�H��7�ղ՘k't�/3j�'����Y�	�:�@�"�j�:4q$q��}Q��O�_�px����:�i��11�؜/q���C¦x���4�����BUnJ��*� C�j,F_��>�!�),a1��@�2������G��DG��}�ʨ�t���lX=�p�J9Ŭ�/tJ����3y>[6��n;�N!)[���[Lj�wS��;�t)�s��p���X�E���;Wv
3��d���.���_�
`����%W�۬�f��M�����j��3xO��qi?P�DjN�����)�ܷˀ�[t&�	]�ڃ�pAܛO���xQ/Dq疙��̍���kuW|/����5�hK�AVg�5k^����q�������}^'	���ƞZ;�u%�t�r"�T���x��J�K	�-�|�A�� zV��,?�_���5��T'�WD]R��,�B-�Kgl\g\bOe�0�yB�<ѽ�
f]��{B93�o sl*6���0�� �5K�0�E�?���2�Y_�ڹ�:^�����es�A7�[�?y�fDB%�����{	%,=
��]@d8�G����������Қ]�481 �Q��J�4.{7�ZRݍ�F�VvO-���Ң�=Ő����N{q��� �j5׮�5#�Ӎ@�۳����È�a��SP����`>�E��������{Z�~(b�����np.&[#-�E4��B(����A�M�W8]R����T~��(���v�h�"W�{���M�d��)*c_Y�8�ʟH�A�t�!�*���AtV����߀����:����k��s`N������"s�b�}���,�.t����!dfB4��$��5(a߶�u�l�ZP��!��&���Mw>���k��[-mC����J5iky��;bHv@��XW����Ƥ>� ��Mc�)y��@Zi|!��I뇨�2�������3%�6 <Tگ���K�}���������xz�޾��Z��S��u½�Z�v*�����{�sǢ���4V�b����^��mг��k���\�{��N�զI��}4��;��խY�WDS����o�w7oQ��,LS�D|@�d(w�$�nSA	��8���+o���k��Ȓ*���AN�n�/y�9-�
�2�J��0��())�{��j|=i�}dWJH��D��y\?p��FAޏ!-�8�$�}��zQ�"��=��Y.�)!:�u[2��z����4�3��h8�!RS`�h�h�P8�X��P���/&Fj� e��}oɞ�������*�Y �y������1h�3y^3k��u�( Fc��}7}��O} �z�'wk�ל����&6d̠�(����V�eaED�x�d�b�$(���z���TG����,�Y@��~��}�r��]r�r�vt��zB�$j[g)
��s{����a��3���3���DNM�Y�	�&tu|�[�0x��m�����5�C���n�k8u�K�-�j�������H���fo�C/���	�d�� ,U�4X�GF��)��P�rN�{�;:�<q���sBz'�<�9~��.����j��]�7(�! �5�j(�]EN*��=f>��w=T��" 0�{�O���NnЩ��d���e���h�59�J̀�;�����쯛g��wl&�9~jn#��0�)^W*���r�i��b��G*'��k��Wl�=�� e�U�x�u���;�f!z�\�lS
�|��G�:_<a�Ԕ��h�<�����������͋�5����4��?�S�yP4/OH�����JtD��n��P�%��.0�C4s=����-ϻ�%��Jt�`h�6^W2JN�S�
¥ը��g�C+9m�mG�>��˲�3�	yOt'۫��ڃ� &%�F6yY�=D,6�l\����-�`&-T�v��Hx4�s=�����	v�iHx}Բ���&�a4�v�%�L��[��Bӆ��1��l��[&����:�H��n���HD�Ql���L$�����,ϒ'M�F��z�f���3��� tb�~��m��m�K��b���r2�.BSA7t����2-����Q��`�|�;a)����F���̗��&��z��.�/����jֲ1�џPB<��ڐX�i�B�c��c��x����r�	��4��Af��p���(� ��X5�=}J֡��k�ߓ�RJ��9w���w'��;�t��պ�|~�v%�uc<	�YӇ�S��V.la(�����lK�O�S�LvYΑ^c���5#DID�zH��B_�8=rf��|�V׹�$�UvRL{�[.�(����&�9ٴ*��,�K�0vV���!x:9�G�BB��gMN�I��Z(�Lc�;?ڜ�Ok�QoGF�:�׸�9�166u|����'�@�r������gJ������9�������H;&HĿ�2�����Vfa�{qkl�~�Ϻ��������7X��u����O��j�i�Mp a��VC��p�Qԓ��DC�2�a��-ʽ,k�n��{����Cq2ӟ<��W|1�vW���Gy��)�G_VU�&�tH�a�u�I��k��	���6i�씮���U+X� ý��F
9A��>�%]1�dT!ϑwr�8@z����K�{�rj�xF�I��5^�垫�J�U9o�?�����(�Zy^�iqH�6z�e�����꺣�`���_��t�6z�眱v;�����vؾ�u)V;�S�3�>��Ƿ0�%5С@n�z���V�߮��D��&v���;jO���|b�C��$�FP�6���q��2�tp�o�5s�̮���Jځ������hY4��b������I|S�E��!���$=�����ZK5׹��{Ʉ��P��~����ɔ�?Ǔ�6/�
uO�K��Rq����R�W�p�Ӗ����rt\�4�qv�d�zhG�����C { ���aIv��W�B/ʃ�yg���X �����x�7��F�p[����"���A�x�3���YI(~g��p�Xb���T�Que+�I�w���N7���N5x%D#��`��[CL5N���4��I�ay����B�y�j:)���!����u��G��-����c|�C$��P�/�