XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��2T��G�8��h��O��ϝt�(8�h��b��)���+<�Pfi��	e��.S�hA�AR��gP5V���9�6���Ká�X���u�e��[�G�VQdO'����u���4P�oX�SI�k�� �\!�!h3��b>^��֭��j���ūJ�3J*�S4���O����A��hs_��h$��M[���9Z2��/)~��:����J�3�$�+fj�S�~����4�<���ّ#���,�E'���$��g_3�O2���c8
��
}����B(u�s�����'���35����-Qek����}��rx�V��`���)m,sEݕ���i�"[U��<�('��4��5��ܳ������>Y������IȲ�DC)ٯ0qXGu,d��yDF���Ԙ)�T
K�Z�v�(��ά�5o}�`r˓��y�A�Hr]���I�27�ðh�jF<�;��F��k�$���ʶ�U`�q!:}t��g���y.k?%e�6��3����Z�m�l�wSZ?�D/�c$%=Rꩰ���%#7����߶�I	��@X�Q�B���0hEz[j�3��/�,Ak��gR��.W5��n����*?�v�p� �!�"�s�AzHXV���C8��9��`��=&EB�P얭`�q+wIǏ�pD�������ђ=�Ϯ���ƍ�L�(SwA�\V��~J֠���V[��8��k��!x5#}yg�������8���Ç����eUB`�XlxVHYEB    fa00    2a40�-�~-I��/$sN�Uي��)�5T=Qg���;\1.��b&��G\��-[�6�h���:�q����Z���Z��p"A ~p�F�K��⬥�S�`���6��]w̚�ɨ�C��3���v��y���'����Ԥ$��07����P�J�oX�T�R����w�<�x��r{S�&�L��Y+��Z��u�	D�C�;�C�)�q#�fa�*R����7�D�+ۜ�V=5�"�|�
A)��������q-7h�.��u��H����׳���ۃ�>��!��e�80_�{�Mv��Zu�����H.�����{���C��^d��5��]�|�mgH)����ֹ���N����XحG�a�Ŗg�J��9��+�[�M|�K�_s���s�˳������$��Em�e�M�a]&�/�L�z���Y��d��Rltf��]����?��k�5P�'�X��
�,w�yьu�+}T6^���5��D1�I�hg#>v�y��O���������ߵY������?���J<��>������#tc����b
��d��Ea��@�B����=�oƃ�*�8�k�E�֣�äy�!�� �����委?�rg�`�P��~(��+b�{`��4���/Q��z����wa�@����˃D��S4���nP��Y�s��	i{�ɬ���i�j��
�a(�]���i-�>I��T�='CCf�+v�T�n�Z淔���(e�L��t�}�U�_��{�S���ča��m�Kж5��Z@��p?�j~�ՌƯ����V"�l�n	v�Q�]-t�B�חS��ףS����2v��O,[��Ԡ�0����"�3�0�چjY�h:'ft����m�N�*��ƥ�&�s;Y6S�e��H�^��r��qY�ݴ�Q���g�ť������^M�������j�c!_� �Z٧�䟪u�y�
�^[��H|�N�m�M����h(Ό������D�zk��/��f�%��@6+&2C�Đ��[��9n���P��|���ت+[�Jr���r��(N9LJ$���F���FтH6�	�;�e�䃪x��8�9�K�R��>&��Y�3�������/�A]c��n���wPp�l{OL�QYRr�ۗD�#����qQ,��r�	ieژ��k�FhЛ8)��V1]Vz�]VTPvz8p�Hz	�+�n�T� ��stq�7���cK���*���a��b肭x�Kę-+i�D��fׂ�C�����I)�ZBL	bt�cl�A�Ho��A�u�N��[ʘ�[��h���E$�|S�8~my�+!�Ay�8LA���9'HT+%�#��MU[�J��?6ˠ����c��� \B�ey��"�����$ew4�G!��vS������:�p��j%��<�PV\-�e��퇒xİ�<'�*�I'�(9��>'�=R�LA�!�@�;^�>V��<��B��"I����/"���Ƞ�N9����X����=)��#��z����f�o����O�c�:��37s�3U���<'v��
WT �����k�[Y<>1!����!\.��V2}Q��-4=��F�N�4�:��*�B�_���)d��k�*Uj)�&��HB��ژ����x�QE-7+~/@��?�r��ӯg<��~4f�rD��ќ� k�O�g0��,�>��]ؤv���@��P�2�Bo�j���<�?���6�/��/Y@�/At#��D�/@cAe'��P��;9��Kf^�fq[ק�:���g�~48��H�܊ ���:E?�g�<�^*� ����[���H	<������_N4�BMw`�?*�౅[�]���'n�m9�� A�yO�Īp ��U4͒$$����,��NY�]�����o-
��������.SM��~Ѩ����K���Zt��ӗn��x1.���M`�1)u�&���r�3����O� ��jn:��)ױ�3�;���8���m���E�Up���4.}���X��e�h�6�鳓qΦq��)���������*E�T��͗�t��ݑ���Y�{��؝D&�=���+�귳S���^̍��C��8��֏bLR ��I�lP������`6:w���,�^��/7\L�.)�@�JY�i��[�^�b㥅�1JQwМt�7ʥ������_�xc�����:.}gA �R'U�7�F2�+�҄�-�Z��$�:Jξ�)7��T%�g^�j�Z��.��F����J-]��J�d7v��Q����լo�ܔ�Z��-':�;rCq�r�
qv^}a|>h��K�ѽ�һ�ܭ�Yw����A�*��\5�^H��G�s<Eв5:B�y��
�F�gc�C�$�1e��C�#e�j��Oա�~��'2ŀ�,�L ��5�l�u:m��ɘw0�t�͓26�(���6���$��rW���1��i����i�i�~�
�g�1e�n��}�m@����n�p��tI�J-�yB�e*��<q������N�������{ā�����H5�������!F�e��?C������Lx-��`��_�c��/ͪ��׌NP~/[��7H�~i�-�����:���r6�oC�o �S�	���\��rᘫ#ߑ��&'m��,�A�U�iy7Q�m�R�Z�qҘצZd8����Q{��i�v��k>�7��f�娩R�� �q��V��b��@�Z��hm��6\�-ܒ�
T}���R��/��h�50�lq���ʒth"���t�%��� ��6.\T�"4��:���L(NK�/Q�8P*(׬Ƥ�EPnd��b��&^-3&�6��=sA�y{���R"CM�:|�Q��Iu� pnS,NcJ��%�=]8��,��$E�����3=2�Wzњy��,h�k`�%t���]��3��N�Nd��$X���u��.��M��V�`.Q�U1�?��R��S�ء	�i���q�6&�������^�8�$J��{\;ƀ"��'"a�HM �lz�t� z���@��x!�ax���H�	c����[r�T��ˎ�yZ�2(�{	���<EU���7ݣa��"�@tȠ�q����b�QY�.����z0;eL�x��.���ј����U�)�?��Il1� �4�9���W3��Y�"�}�u����B��a�3co:>7�Y�&�9}S�����4 Y!�'�"!��	IF_��;�
��=��維?�jYH����,>���]�qy��Z%),�#��N(BK�����z=��{���vc�9Zl���kv��J��fD�R���-��B�mu�N��y�t�{�T%[�8��A,�7��?��Bb�̝mZ�5߽O���:�a�O�-qR���V����n; x�tl?�j9M��?�Z�,Ƿ�Y1Zv{%Q~����������'s�|3RB~��ie�g��q���DI�C����՘��y.�;ض��T��v�����^�����\�W�Ɉ'Q��1��W�r+�� ����[ň-��ٲ��dD��Qk3��w������|���_���߀Iٯ⣭x������O���4!A9W$\@'� u7t���:�{3�rސ����a�����98���L���� (��\]1M�ML�V�kg��ѬQ���/�M��a�2�uYX!W�����L{-�;6DG) Ch��5����DSa�sg�X<YV:,C�_���)����#DM~�����sO��x^�{q�QՓ���.W���^�+cjT�6���>Bɡ7F܋:;��|����g�����͠��'W��<�!1�y|/���繦"��ݴ�(M�؊YB�QQY���
�0j5�N���"	��p� 
5Y����"`]���q��t�)��R��Dg�PgjX1C����l�T�'�"0�B�>����uN�ډVO�V=�h.��揈����B����v���-�ڭ���=�1d��8���/7����\ǻ��vl��m��6Q��?���&AO�+�g�a�!srT�^��b��eA^y�4��ٯ��^��7��Ea�6[�;��#v.�i���sSX�MO2��~qyk�P�-�m�$���W�@��<Q9�1pN7ԅXB���pӣ ։?u������*ī�q��!��W���o#�d1ωho5/ P\�Y:^�W��>�\�~Z�Nkl�m��W�޶t}�Zf}o��u���z�q��'�s����~�`#9�<�鳰.�}�!v�	��`
˫�C�[�[Í��!���|�0'�i`���'1)�Pn4�?s�g�j���4\!۴��\x�����KyJYA��\��#�[F�/}0���h�Caq��,�ʹ�೚	��Bl����a�eq�@�o�Gv��Z���fc�]��H���n���ʷ�,L*�i29_b
�����y	X��������<ܚ1P�^�0��1 �K]eB� �_L{�&����?	���7��Z�E�1�w�D��m���;�M����₰��k� V�0�d߷����M��4��?��{ｰQ�vV3�;1З����t�)	{mq�Y�� ��d��̊�作w�١E�n�_�93in�.-E��s �ذ�=dC�y���p��xc2�[��A�h٘e~�W�-�h�^:R����E,) ����9o�wҮf���<�����L��aq Y��2�J�`�.]0:}�ڸ�e��
�kp�!�����)��	�� \oq/�jG*'��%5�r}�Ԉ��F?m#��"�E�����o��h�	��_�5����<)��r$��c#v�2
Z�U�6P�pY\�Ҝ5��{�#��\��Ѕ���	nA�em&a�&mb3�֐r���ۊ�Pg�]�����^U�o9�H������0,y��d�`E�oT$�t��ٚz`� �x�z�f.�Aȟ$דh�o�Uv`�-�㌁c����vŉ�"T�2��� *0k���#��F���BN�"u�-;�jyS�$!P�7x+���{`��@��g���5�$fG,=s���d�]�n�N,��)/����cz��`r�|.��ʁ�U6H��7u��JN��	���t� 9e���V�7�a��n��Nnv�īƑ�����x��|3 ����,�j}����R�=��O�(�δ��;��4E�mf���۾�h�K��t=ad[�a�I�#�ytν�G�W5��V�������":�˦3��+): �Ck�B	<����Y$/y�	��W�V�z���M�������v�l���P ��x~f��x�S��Z"a�Ir8�a�v���֨�����������%b�2���2�R[bp�~����V��IЏ�ۤz���~�����ԯ�
[���"�-��x����!��n��Uo��߸Q)��"���s�y��7Lٽ����L$>A1,?����|��7��Sl��F<u�3��gnG��Hڡ��1���P�:�%�m�~v1z}�E[��:�G(�W8T���ua�4�u(��'�|�S����z�J�Yt��>�� ݲ��G?1��?]��6@hE��{�:N���hIω�+#����Oc����i�5�����8�#�}>�e��褲`��'��I(r`Z����n]�?%�b�}H>������K�=Mi@�Ҍ���ZsrCU[�?����B�b�xlHTcL�Mݪ0�޸��ľ!����x��F�=Z��#�싼ş��W�;&�M�j��Ah��0i���!�h��>��o���3��[�n�H[�.�,�*ت�҂옏DR<��{1ޘ.c#xӓ�<s���X��BI�B�,�e������8c^壘�訉O��gc�G>lW��X^���Ut;���0f��"sl潞��樆�g�`�qA�_-.�K��ƍ�Q��C*�*e�;K �c-�/�d��YMi��2I��Û�'y�ϝn��R�U���BeX+kT��
�ſu�@��h�m����k�	�X[-�wMX�J^����{�X��E
w-P��LY�=t����t��O(2�'�{&%��ӝ-���:�� 5�.�ҀC����jj�S�Y��O�������b�.����/�‌��1��b�F!�k9�������T��*��F��䜴�ߍ�s��9Fp�q�6�Ԣ�B�aHX��e�s�&�7��l����)��R�.Ŭ���I�Z��H�]���c�drjF>�h�y�'
\2ʬ?
��&8���s$t>�ܺH$W��W�8�3�w�!�I�a���w�\��!`}$z-�ȭ�����A�b��~u�=d�=M)��8 �*����-r��Z;�ѩ�N�S��t���X�M$h鈞@2d��	������ۨ_,�R��3zI����L�b+�|T�n	ɽ��>�o�$% i���U�0u���o���]�܍�R~cg�B.Ѽ��Z�6�Z�yu0�Y�,��w�#���	�`��ˍn��X�������m	q`��G��B����S3fb�ܝ�F��2o�Lo"9��@E����پ~�'.:�4��������At8&���Qd�#F�z�=e�r��N�\�TG��l��)aɻ�o�����?u�~�,>�AQ�rخt�&��ir�7[��W�T��v��H���� "Uƽ[쪱����' �hV��U�
�u�9/�_��U�s�ɔku*��;�᷂�Ҍ�U�k�c�h%�<HJh/��i�w�[�$c
�T����e�^��@`��f�Ȇ���ꟁ؉��XV�N�V��k��E��T���&:��Qָ�6�[̱�bCs���Y��[AvnA0qC��!J���L�!2��'�d�/�ܠIͨ.��q���w �����;��hZy��=RQ/�-a\�]����,��5Y0��J��잫N0[��f��.����� �$_;�i:O"YYr3�gOc<����F���/ F�s]���M�O�ȳyژ�Ϛ��DI�8]�6�ʎ�O�3�{+N-I+j���A�&�<�C��@���;�4�5��27���&�ӊf=n�~�n� �]!��m3=�5��S�6���*���H�^j�n�H��p���|�մ�C��G���Z�s����V����赣|Z�^r�S�D��/d1�	`���(�c��b8�}��M:6�"�.�.��独�"_�w<����"��+��]��Q����]VI�
�ʀ���(e�ᅑsHD��੥��JY�m1W�N˻	P
��$J0y�@��Ni�;Jѩ��K�,2��ⲹeH�Ks�NHN/w߭	�=X�7M����N_n#u�D�-����?*�Ȭ�Qݔ;�ʗ��Y*+��������H�\��4&�����q0J���ߨ�ڷ�:�v#\C��}U[����߅2�D�]�b�]"
�A/sw��9�tv��0�u�b�x�[��˴�7⨬���y�1�ʆM�fc�ں�R�!^�N4%thW�sV���i1�A�{I��e�Q�룛Yh�|)=�B� �<��� d��q��2�B�F�<�yA��^X����Ce�U���\��}k*O����<��%�Y����r�U��xڶ�}ʂ�������ڷ�*�@�E�\��RY	�W��Jc�Һ��)c�z�@p�*��f�k�Ϋx��(NS�HB�5cr��:�����k�qw�2=�B�'�1-;�N��L��hW�w<�S�_�.�`�$��Y�P+�\�:C�J���Plu�G!>w���]N��A"���;�p�׃X�ۇ*���E8�m�3���720��p�/ì7o�c}k��O�`�00�#U�!G�]���g������q�%ט�I��Z�{�. ⫧͗��a5��8ߪ�<^g?�	�p�����2��2�R��J���}j���^��U����;���8�4�\�FD�GI��<�a�wz�hp��E�^u̯��d�-T�
]$��g�츝Cx�_��a�,P��Fn��}nB�ɫP��/yz�����ďN���f6��Xe��D��oS�.E�rۗy�`<:��%˟-C�q���s�A��
���gvf��:W��Rx����sD��E�ബW(Y�Zj!j���{�7p�7���&z���� �3(}�P�Y�	�Q�����;�`���g
���Fп 퇫�������b|�J���������]�&�B���zZC����`�z��˩"�m4�N]Ũx=��:����=���F	V:a��6_��V'�ř���@q�,����6�E��������{���!3���ʣe�<I���v�Bh��� }�ہ��·���~D����"g7�=w�hvv�}�آ>��V��Lz�hr�pU��a@g�6�ws��gndO�gOy�E�eԤE�ճ�　p}3���S��f ��BB�O$6����f7C[l��8v@�!�Ɇh��a��U�N�Ԛ�R �BaiM�T���}(�d�@��]�����뇝�G6Dsf���ʦ���?J��h��4�G�'-����<X�}��j���`���ó���{P��vlY�8�C���� ��Q�!��g��is�^�Ԥu�:Ǚ�f�A	|�L�wii�����ؑ���c��SR��nH��׺�Z��m+�����TT0q�*���.M�ۑ����y��c����� "Jm�M
�뇻�Dζ�Wt27���#��%����+,.n���,�;\р���*<$iY���:J����/n�,j�tC��'�L�/7�Q6�n�ΰ�`<�!��i�����#"�&�^��������ω8�/-.̰��ҝ����И}Z��ئ4�2����d�U�|%J(ں������+H5��s a�D'$�V,�C�%}V4�u�����~mf�p�ʇ;���c���љ�����$h�)�ޘ��ې�ԕ��\�y��������P,j��O�s��wVH
)c���e�r���e�}������:��J��,ǈ�����lFݛ!��+Ax-�@OW�h4ʚ���FDO���z��Y���|=(,�rV\
/Hp�[��\
���E���i~��'�3.���=~ �O��AS�x?1/��ی�8�\�|��@�&h����ԄH�����S�+�w3\��UƱ�J�r9��J�G41��2��2���*]��5ld��g�����F3a��Ԫ�M��Z�5.�c�>m�?>X/�.X�1�-�_�h
�n+<J���D�z�u���q&�����*^���Y�ծ����~�#��"M@2M��w���iӾRP1���Z�3�����c_��\�{�p�-|ex�����+~�U:9ɲ_ۻ�ӊp����?D>b�ߛ@�<ݚ��*�D�#�����U�;��v_�b�P���@��PEƄYJ�I�D��&����/�a�P�Q#mս]8�e��ԥ�+��a�(*���NG�2����lP}3ۃ`�h��M�9�Y���y��r�73ʀ^���A<˧Y��j�x�(|+������ʩ��{����F�Nb�(���'úb˷�W��d6}���7߳��Zd�fL��\�lč�;-�}"���@�K��¸��F7t�c(n[7���W�2���C]
�G/a�z�S;�}�=?rZ/Ћ�r�$ڱ��Gx�տ�3 ��Om%�H��b����](_8����>M�`�i�(��$�*��0�!�Y*N� �(%{�[�P�B���ݼ�Kn`��ß���@��C�9A���ԻP_���gQ��o�l���F��n�~Z�ׅ��l?��-;����EVڭ��3�Ӽ�8�xdƇWj34��7�g�t�+����.�IiN0��c�����7�S�鲥PD���Ⱦ��c�����K���H9�x�*��ߪVc��*���ا�/��p4
�Lt���5D��<Bg�,o�*�,.�	0�������'���˴����c�>�2��S�ں��:���SҐ9t."zH��#$.������e��=���1�l�uɭ?셖���J`��-�
>]4�	���q\��TR�#��Gƫ?�5����D����&Z/�Kf�t���D��� ��Fw#����IO:���v����ս�
�y�8�$lI�0�y��g.�ıl�f�Dn��`h�$�{���R<o� �����kUq6�F��X���u��sd�+m�z����Ƈ ���ӫ�ꪝ�vt����E\2�d��"o^#4T�mك��� �r��u������@�gӶ�zt{;�����\w�����4�����D�Z5>�=�3���l����/����E"�� ����6%���Ch�We��Q{Y��6�	O{��N
̲ɼ�gO�4(~�����'<��}/5�q�9�3u�����]��TIWZ��1�7_R�
O��b9� ��Q�T�ԛ�x���v��<�G�Ǘ�1ˋflh1_j	^|�U�-�E����L�^��� _rd��{f�gv감X�C$��M�.�v�X�v�կẏUѿ��b�����u�*mm�-в��p,����i�x��eŐ5U���``}�: ��lȕZ�ȶ��c��Av�2ϊ�=���;B�)�Q2�"�syD�{L�XlxVHYEB    fa00     8e0�����������{v�5����8������]��ac� ��d�8F���9+�*�!u)z�wE������3�0k�@\gz���Q(T���񄗎>ʼ��|�8����4�����yF��J��M>y?/��T-��������}�h7���a��/��*Z627��ȳ��)_����aas7�3����,Y.涺���>��M��̧R�����F�˛�o�0:�zUFR!R��[�KZ3YISa�=��R���a2՚M��~�N�	i�)��n:��[;"(��&C�!�։G����>����'�����r����Xb��Vo��p��Ȣߋ2�G��;luS�J��ؓ}��	{�y�ڞ�$M���!�oH^���5;�N�NC�����c�`1��������O�Cc���'�`2ơ��8[1E��}fq��7���Z6a�#M�U�|-;H7g��]XmV���o������B0{����ъ`���r7{�[�ġ^�*���x ���&p;/�P�]=���rt�Z.���.|4�.C^˔��4Lp��b܋�T.r�u��L3���4��P�JY��Av(�n��f�Tt��
���ݖ7џ~	�Sa�d����`���.���I��z`XS�@�;�#�e��:��*�M.V�A`U�w�-d�t7������s.�����W�~)�.M�W�p�˖�X�B�lbV��1�8öv��ۑ��z(����6;D�E}�9�Ƿok��hC��~�?y��,E~HN�WCA�K�L&ԔM���6z���+�3����B�Ke�@z��Qml�b{y�!h"vao�A��M�V��(�*ؑ�gy�O�{�3V�B�z��\�[�=y�ѵ���zS�'��Q��V>_�e����N��T�]^��a����`^�Y ��w�)-�����Q&oD���x7T�w��i���c���3r��@B[!��=�3G�Lj��[�geD{�Y�"�ӥ��/F��i����lt�V���Kpg�mĂ��4�:0�����.+���7�X�8-x�9��p߉F��3�+������hA��3���@u��<<W�XLO�p�2y�&�C	]�[+��ؒ����w�G�U4�
�5y�2��{i��>�����{���>�*�����E��bש;�X�/}��0���ژ˝�%�U1�V(��c�/�0h����� 1ݖ�D�s��U���Գ�2+�f���D����F��,Fa)6��9 �Q�q/���?nD��ߙ4/_�z�����T���ur8�X؞?�F��$���R
st;c��Bs��Y�B7z0	%'@�*��%��uyư�%�;�1��Z�QR[Qb��2���ӚxE�bյ2CC&�J�����;��v�<ۅ�}�}��+B�����r���.|h=v*N3y�a��_`�� �_0�9BmV�+xh��
���)��i���]�XG�$|�'�|"����S�)}
�FP�		q\A�t3�I�-�%)��(	�.�� q��9�S}		h�I��-椎�g�Y�g��X�� �{aÁ��U� ���`D�a���$��:�[c�����/�;�=���,���r�Y�. �u=i:ln֯3�/_�Ų���g��?���'х���֤��\���6Ǵ��°s�ĲтhY��L�Lu�n��xxf���Q��!I@���\�eQm-��Z~7K�r�0���x�!'��Z��\N_����/��u$��Q��Xߞ�V5U�%�Î��z�k�%w���]RS��aZ�� :�yl�Z��3�zE��3�}},H�#p��+�n\M2��ױ��l��P)4�Tf[/��a�b�ТZi(]5a`��:ad��6��r��G�m&ua]�G��&*yA��k���ٙR��]h:�T�x/�
�[� ��1Pw3;e^�j�ٗ� ѕ��졆Bܔt�q�Ÿd�u%����׳�c_�C��D�������1�P�C���=��a�d^�˸�N	��mA �+
�׆�>����w�N*1T@i��K�V�Hh���|���柾�������Q�z��Nu^3�)�Ɩ�9��+�V{Z����6$bhY~�u�Φo�κ6�y�}�iΏ�{M̴Zu�IJ�1}~lC��D�(������N1w5���H#Iz&�dL�Z?�|�!��l���<P��4�6�@+�g�	"݀��[�d}j�twXlxVHYEB    fa00    1110�7[� ��3Ȫ���WIv������o��c]5�w����&��뤍�*�)��n!�ndR������&�C^T��
D42�[�#I� ��G�b�+z�T��O�Aӊ�mK�im�T��v��~�㭦�	�uܘ��p����/��|�r �V�O�a�%y�j
ɳ�=5)����9jrtL�V�Gi=ҙ���e-|A�IN{�`�?!�%������ H��`/ܹ���U"?u��^�_DT@JV�q=���d��8�6틫�1c�ޭ���2��C�-��c��4S�'���R��q��*��Y0�{m�RwGl�����a#�ԥJ������^2�F�D18���b�,�ن���˙�}�Ռ���.j�[VF��j��<�#�yF�S���>A1/(X��@�TBA<�hjͳt���ﴦ8�>ҕ᫓J����JhC�4U:���	NI��k�G��E��0?l�OV]]<ħQC(��Qj��r1�I&1W�Zń����7��4]�/2���nC�e�}j&��b.�@��f��X���6�)�$0ۖ�0�߹�-B�=kd�hc�;GɓT��v�������VSH>k{= ��fJ��X�W1�5+�6���E͓���M�拫�D6�w&�↞5|�#�-I �6Lk��eX���b�P9��O���,�A��!jA��v�\�+���K;t㔏̅Jk�3$/��a�&�3dj�a����xٚ'H�`,�z�V�08��D�Iִ݊SeP��n��CI1غݗ�*���M�B���ab2�X	�N����kR�{���㙠�4C��a ����fڦ	/qw$=D%~��+X{'�}�l���S��-��'�w�C�ͼ�i�W	eau�!i�r/a�q�D`��-λwk�0]�;"�.x�ux���R�z��2Q�`���bi�V�h$��8��G��I��܀��s�-R9m��m3X��)ұ*�a������]��lWQ���^�P�)������n�uW���w Y�0S����
k"��^7a�ɥ	�Tmג,��:!C�0�oKЃfmfbM{�w �E����ٛ�&z���jw��/5Դ�e��/�^���,<�n��؄�����.x�c��g��+���A/�S�87b���ç�r��&A1o�ⱦ},=r�P���	tƪ�$��T��/Љ(%�1�(�a�ݿ��!�ձh`�ʷ�-��9�j���3tfIj�qn0�b��&�8�藊)��ǑS�ˢ�s�#W�k�E
S�L?���@�ݴ,'�@tm���_�׭9� �z��k�C��F���x�,�["X���u�0w�$d{N�r�E��g �	�7_���y��P�P=mk-;���)|[�d)�{��ϟ�����Xhv5�I��BQċ�cy�K���v"P����S#��E	X�4Tet��N%��̹]�b��>\۷�j�dkA��¥��F.%�

�D��B�~Ď�,�3t�f �4�a���3uH�o�_�B���a8R_.h�oh��z�==����,�6O�����'�v�ĺt��˕?��a{��Xr��ln^�D��0$בX�g�ȁ�.�j�D2;��������#yMS��Xw�ۏ d��l�k�/�w�<��Z�57��;W�]�3�֬�V��x��;jJ��^����r�?̆�װM�*9�� � oa"��� V�����Zco������9dג����bwm�:�e�P�)F�H�1�k����l�ocf<����>z�V�=T? �,�b�����S|O�-|�pY.��G]�N���t��⚲�,�B� ����ʞ�����x�T�����������-A)��l]��Ό�!�F]�7!X*hO�s�J�U��t�!q�v�}�/o�r�HM�f?�Z�6�I��[V�{����W��9���WF+T �B�SQ�>�Afڒ)?�\�����VG;p�:䞝+�ɛ_�����-;�,r2��C�}q����x�ºH�������c�7zޞ����G�m�A�U��V�n��ۀ�'\�\s֯���U�]�^��P���n��: Հc�f:��l���o2(�R�~yv1� ���>	�!IG�:�Ę����S���(U.V�#�@a�̄��"⺩�TP;r$���H�'��l���E�\��(������� ,F$cv�A�z��}ؚ�<+��Rq���In+?�v>�.6���y}	�d7�K3���˽"ޡ���D�ZҐZR�����'�N�
�*��M���%5��J�pw���wӤ/�@8z�Հ�k�D.,����H�V�Q��)�c�#��>��	�'�K�����pf�+����z���T|�T���a���˝���y-M���̱���Cr���ڝ�\HQ���:���?�C��`8a��1q�wu ��B�N�E{\�)�Ύ��q=�٣`�D�6�4�C�;�ل䀝
���ך���8p�v��Q��֙���=�כ��=�0�n/H��q��P���l��9x*�`��Ov����X-]�/p�:%%�2�	Hϸ�	�dB��1�Dw�/b��r���fəR��k 9Ҩ����(��J����ۡ�gB����"�Ho/5�9�������O��I��{5�������Q1�`X�Uޒ�Nm�C^�55v�6�]9���?(�*%��q�t���g7D�]�_�FgY��LN���$�h���3j	~��آ�3�#:���#4�I�\_&�o�:j\
���6I���'�����k�+���� JKav��i�_�22�.��d������ ����?\6�W@��⦾�.H2�o(��r���N��b����D�䌋�V����idQ���	,o8��m�H�_'��#g�=�����q��
�����&���[2o^�g���o �~��Q����Re�g� w���[2�� � �=Ѕ�n �o��ч[����R׺�c��5�ꓮ��.m���sn��G�l~��'��jv���g�X,��Q5���X~w}.��xW��t��)P?<a;J�1fa��e@
{��і3AH���ş+!�n�B�� s
g<�C	Z���
� F&�ك��0��x����)0;�j�E�긥��~l(�'8����P�@��Q�W����O\��$��֠u6�'�W��k���?:U����E��B�/p��Z���_b��߱��9���5̅i� F2U�1�g8MP��0~���x�誠�`�t	[�`�W�@�zzк�悭a�?Ej�^v��OIzV�7��mk��N�7D2X���}�|��%�]b`L�] �5S�������{��R�<.��}���UփUTh�&��;;��=�g��\^ۼ9��t2��)D�h���z�`ʝ�`�0IȂ��H�|����+���H\."2���n�vS��n��i|���C�P��=�>���Q�Qv���}
)c ��OeJe,�=�0�@�8Lj JwLGd�:�~�.0Iǁ�c�]M�'�v�%�'>�S��[���ܵ[�8��hĆ����a�_���ʋ�5���ڌ8J��l�$n��=��� ٣���ڕH���Cȅ�H)'nnݱe�#!ǠF�ː̾:R!"�Ӽ/\�{�[��܎�3�ݔ��~cf�7��h?w�G���r�ļ^ps�7hk�0v��}���������8�k��x\��7cG�z���UBΙ����%�I*μ};K.�-��ǜ��E��b!}�i�I�����c[�|��?�:�m�պ�>��hc�bu�����>�-���Tp-:Q��U��M�'Y�T��J�7��H*�β7m㸸$��~��Τ���s28�L ������W����.�k*dB%#�������W.�u+����n$���&_yr��ڞMm��Q�Y� )��L-R���t��Ơ����k��������g��'�p�Ġw�E�K���m���^��{}��?KX2�{ ytE�A��Ȩ*�Q�)��'=�c���Yg��Z�~��0�4�JƮ;����6�oN�N����>�f#+��n�w���mOR8�A���0O�g�'X�|x��F���6G٬�e�)|����W��`py+��1����>w� �'	u^�(�[F4�l(]�[� [Ե bc������ݹa�
��(�0Y�	Qٕi�}Y��كhξi�}C��K�N�l��Ǿ�9˯-�3]���#�XOLhP��1�_�ӑܙ ��4j+b�"c+<�����,���KJ��������kh~<�ŗ(��)̋侖l[�A�XlxVHYEB    fa00     ca0�4�մ��y��ƹ�ؒ3�[@��C�;�&��2~6N���!1����rA�������[�B(uy�վ�X
p(u#I�<K����uoo���r�>��}����e(i[O!ʌ�ۙ]y����K�b#�C�{�}���Ǝl��P P�j��K�#�����t�+3G�hlѥt��^����-�@SC)_v��7qg��؇�e#H��E�7��C2�����Yӱ���>��1���X��SQJ��0F+��dT��#ĳ�oa�I7�떹B`_B�X�f����XpT�O���'6��,\|�* �,�)�����9�]N� 4s_��Ã��,�����ZX��Ҷ���ա�[�,�3;���s�@G%p
�#n@�P�7��6L)n��Å�b΅��Xtөi'��5��HcL�M�ӽ���Vʅ�����I�F=��������.$��n� %Y�m9��l��ǈ��oz���e�A,t��Y�B��T;�@��}\��کN[6�l�� DM^��X�|��kw��f{X�͝
 ቉H��v��5Q�;&-�K GS�fGP/��f��3$��b�R��2��hӵ���O�����C���eS�M)cێ�i��,��I�7S\�\��3�Q����:P�*@�SPp(�?���ݙ_4u4�g�W3x<�¼��d׭ݛ����Y�-x�����A�It��<Q���C虱U�j�,�S1�T�1�\k�;���/I�$I7����i��@EQx�����!}�����(��0�+X(�YH��ͣ���=T��>Um5v��+�U�[�g��G|U`�Ѫ�ݳb�=(�j��*'����J}���>��oY2��:ʏr/����a�4�.��p��jk��c�縉L�$^�H^u��+ �}s��{>�z���u<����=}��=�h��\�4ዉd���	�J��ѿ�a��E��_�4�پ��4�4m��I�yW�t_4�u{�asQa��O"���Ǿ>�Q�=�V�(ވn�d�P��W���{c0���Y�T�e��cM�2�D �|7�wYf;�w�{u|���dg�`&9K�$1�¾0�cz��{tZcV�7��&'��غ�G���UR�a�VDP���P��eK��i��0a}��ve`i0�]J=�@�X�ΈZ�C7����}���wM��=��}���ͺݹ��D�� (�k>�M�B}r|Z�����{��V�����'��rA,Mq��A��D��N	�W�Y�R��\��N�	��T=5�����+���B;��׍�iI�x3�7Y����#�/gG#�K�%��؞����O�8�-	�y�r��Υ?�n�"����ж4��� �Q\����h��u��"T0~��XP2���,�"�De�K8z���^�<�q�����/E{:��ݬ�k���q0��F��Ʀz6q�o�K)��C�a_Nn����X$F�7���ƙ��6(휈��s�Z���7���b�s�K����}���w��=�0��B�x�w�)���?��du@q"�/`�קp�Z������W��q��l����k��{�U��F�2tZ����&@M6�VT��d�7��ꁠ���9��ڌ��P�����+�vNw�?Ƴ�c	z�!�	�O�9�xu�^8c����Ce�rp�.wf�?})�~i1D^+qE�$��\�a���OT�9j���sg�{b%��O�R^9#�5�D��Ԓu[��Xڧ�Sa�����9�v�$�i��o�����H��!��қU�=�`�Ωld�/��C~[�:�Lc���me��NZ@������'��=)�WЙ�~L��:�׸�!�쨤�J��l�����&�W6o�&s��jw �[e��(�&�]���0�������΅
�ܔ��Q_�1ɘnj�Q�+L� ��'';��Y�Aj2�Ej'{�R�h"M��Xtcb��(��L3.� ��6�����[5-��6��w��ec���u�4�C���
�w�-6�kd��m��P�O���t�8�N�m���Č̂�n5�*�������(-KI�y(E�d\�5,�\6*��b�\�G�.��F�}T��֏T4F�v1f~�������������ٛG�7���=<@VG���,�����n��f
�U/ܥC"�q�t���(��,�3V��1q��ze��F�%tpvs���*o~����~p�%��`W���j��j/Fo ���&P3��p)��s˸|H�ʿ:�s"�qy�h"~.F?G|��7���fh7��"S6���!T5�/t�"�'����ǻ�{�}�+�q�)���p��m]�[�{��X����*����wA�C���6=�!-k/5��@�&�%��A���u� ��ڗ�T�JD�m�qߍ�m��8�0����|����'�̑�gw�v�F߶ �	������풁U��T��؂3Up$_�e�1��7{��}�H
��Z��µ�q�ΕSm��<}����[��LP��!��Ut^�z���{s�tmj,�(ŏo#a�>��2ߛK+�؀6��Q[g��h�N�/��`��A&#��ܲ��# `�3�kL�j.��[����Z_�_��pP���B&����s�.�JO��u�Ʊ�q�����q��*���g���w`�5�E-�|1z���H��TSL��Y��'�C�5 �?�G��������%O��Y1L�����X��,hEp^�ʧپ'�@~LU��J ��#I4�s1�`�d֚$gS�ؿ���΅Xh}��|��W�P�6��>QǱ������'�1��\6R
{,���rC3Ɠ�W@r6�QS��HvG�oo�)�h�#Aa X�p&1�^�=M�>};Tj���l�N������ 8]��op�s����8i�1@7n_�AFX�M�A�fM��R�T��[?]R�`�XJ�Q�E&X8�n��Q�o\=�E5@A��Z�߄�_�W���fҥE�e��Z�N��l������Lo-(_֪���� ��{��׋���{����A3�hRk�z��G�}xKʋ�	A,&ֽefn�|��g�������Y>�y|����Ɵ��寤�^$�yPF��817M� ��iۛ����B����T�g�O�68���16��ʤܞ:��U	��p���8�)��G@?p)X��w�qB7�߹�%�]�+XlxVHYEB    fa00     3f0 Q����EF6�y�[��2a��$�X��(�+/5�����VW6���l���2�W���3#��+�G��O�V�8�"�-�H�lwz@Ь��a����V�$���\b�T��S����B���1ˀ���5x\S�ߢ�]&�����rKP��~K����\�]O��̷�Y�P+�����P�����E����f��jAx�,A�DV%�Y-C N.]=ߋ���ʆ��K�⍶3
vPܾ�/L�|T���(�'��V�D;5}o�e�!�2N������7Q�u�B�4SR��A���a�8#��&�������	�m|�9��f���\n_r�=��ν�\3O�������D����}��}Ӥy>�X��iq�DGߚ�$a�V�N��u3��V��x��b��M"�<t���$��~��#w��%�帗~[����M$�%�df� 5o��~J=Q�o�|xj�؉�������yNt8�乆�/z�8�A�ca�;s�:�|�Ǔ�%�-϶�ur����?G�.j��8�i38m�b�.�H|ɻ�\�<G��:gQ����Ƴ�ܮb&���y�u�ʴ�"����zN0��"�:3?j�Cw8�#¿ڨR�7��q�r��>�D��*lg�]�ӵ�)&\捱���]���b���YA��:WD����/M�S��(қ�^�����0�5qryG��^��zr�ѣ�C3�����;f���Լ�@C��9ǁ�Z#������uV�R7�%��@S�gZ�,C��9�'.-Ɔ9'�D�k�|�x)!7GRJA�������4��z�`i�?�0H|K%��/�i�	�l+A�����G�I��ꉃE�'b>I:'�^*?�TL�%ABFZ g�=O{ZVT5�P��;5�vR���(6̂.HA�C�Ӑx �X�����}�����:�	�)��v��:F��Ha�}�;MO���wn���k���O����ӂ�'>W���:ӗXlxVHYEB    8096     b20���=#�f����u��xp���|�t�M��*s˙9CH���� 5�+t�&Y�P���<`�mXH�om��7P�,C~(��*b��00B�Te��1��'�{��^H���.s�t����I�P]�=���=o�J��S__e��f�q��q� 1pC�0��i�݊ec,Q Iw�3�n�a��k�pi��6`>��PQ���
����Y>�q����x�d,uH�	�9�y	�_ɮ�����n�d8��0�\1}�Zԉ��_g��L�!��_��m>b&�����~�� ����'��[`��po5�8�=���)�(�8)Aб�_?�\ӝ�<�>��Zm��� &f�'j��!��1�6?^ O����L ���<m�y�K�x���1���V)�%��y�8>�#�b�l�o���#�^S�8H�H
��#l�5�<
��F��!���v��p��h�>�[�.o�<������b4�3/P ���w��?
�H�\R���S�rcј펈�p������Ҷ@(�y[�fW�6l����8��S ���E.>C���k���9ݳ��������.b�:Z�^��� �Q8�:��~���@~=�,���۳o�1��)->:�m�,�bTnQ���Ӑ+p�1 g��<^_Ӛ�j)[���$ո~��J��9����:��q+��0�e��S�#=Q�*�
�����I!���c]\�����R[��|n@n��Us_�;qU�D�S*8�KR��K�֖�e��*O��o�ٓ�ۓP���y�1���:���U�K�%0g0h���%����/��A�[���Rv�A�m��M ��L�[㔍�h v��#��̦�*U������[�̦��*l�-)�Wc��>xj���m}�yܧ�(]�I��{"�)Cx�s���[�ĮFE����8�:��BY�n�N�$�(��x�x¡�kΈ��L���	�T)��� 1�M�ܜ1A�.EV,}/g������um����ڟ�G�]/X��܈/Ծ>;�4�*W+G�)[�k>:J譿g8���2g�XeN��A-���D��-Y��g���J�32�Th�TaZ.��(�� �8"����i�5aM�BMUl��w��K����G�&�^n~�S�1���aY��zӉS�԰��ÔF�_��)e���\1X �ʀ��';iT1t�2�����A��x+��^{9���%6�E��X�یcl�!U
�2q��p��W�(�D,3����dV=
�D���kI��Vm�ײ�@Kp�&������6�`�(���3���X�.[7���{+VHu��E/�s��,���2撝k��_��sa3�3�)��|r��v �R�.�E��;\k��<����g`���l�d��f�g�l+ġw�Z�+�Է��+��)Z��ԚaA>IV���J�E�q᫈������)�bҿ/;?�̘	�c��x�	�X�i%Wx�x����g�{f�NYzAr��0�@GJ�u�1�dY�$�o�s���2�U�3�4+�cx(aS���vk'�8Q����K����f2w�-�6��˅.�3>��3A]�Y�B�_%�?$B�p�MIU����۵(y�S�tn�,���^�*�e�n�猽Ĩ�s^)kYI���l4ݼ�ڏnB7��a[��>rG7g�7iQ�iÕu+S!�MՏ>�������n}�*J�G{���WOH�đ0�h}�N�du�m���5ݬ���,V��cN��TSqX'C��BiU,��X_7{��9q0>l�^h��n(�6�w$�W�߂6{�@���\lo���E�B
B�HP��4i��gB�vd�
���
~05��:h�b����XCW]t�Cb�<mCy�6�mY��h�V�	��j☆+7� �$���n���-��\
BG+�F�����x|}�9�6"��z�o.[5�ݠ�����ǜk�obqS���~�ǡ�aF�P�'�}�^�[7����Q�&bY����0�A���!���!-kWj��F�UXx;�U�GG�*��(~����ෞp����F�͆�A�Q-2��՜�T������w4�8AvcG����>:���d�ʞ�Pu+!H�.T�X�������No
<���i�����
b��L���:���?���~-��#)}�Z��	����oE�/oh���U>xF<ə��Ŵ���(*"f���Զre\[�Dxb��z �������?�����.�~CW�&c��O�Y�t@�(�������b���5�v�<}��������T�W�q1�i���7&[���L���`�tӓ
%
份�9B-62ӺΨ.2ԡ> ;�L�b_/�������������_�JP{�˹PU|�`���:eY���s<Q�� ({d���F32V� zT���1R	��5���X��� 3L����%} �a+����M��#f�o�?&~O�}�Y@h��2���(�.���n�SK�3�{tb�ײ����Z4�t�7`.�r?(��P�O ��!`�-�5��;iW]���gUs�)P���3j�D�#a��gx�@�]�(Xm�nZ��xQ�~쟇�f	�yhS�Wh4�ð�,VI���/r�XG�l��A��M�K>^�@�#�ݑo�l	�Vo����0��p���ۍXxԾF�F;���d��ɭ n�W�[N��t�V��&S�LLYYTA�-3�xq�������`+/�[���ih#�Ǚ���޸x�O��^�A�&�����.X}�#[���z���.B'W���f��$�t�#�U