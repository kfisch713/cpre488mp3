XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���㥂m1�ᆬ�����\�:�Qt���+� �e�K��v�bvʞD��pߺ�MW�-[RH�1v��$���#%��5�z!$yJ�K�S�r�%+��2({dk�����o�!�y: ��Cw��`s[o����P�y���$�c��O�_�]���Y�)<JB�`kO��JU�@�P�\� �ӥC���!n �)����
�<�*�:�����`�aԦ�ӫ�r�]��;bص�����H���q�1��H|��8=@����-8K�֞Z��vif�ՠLZ���6rGb�+���&�2
�l4��I��F���_�HZ�z$ܟ�+6���S��f�-r9���}�Zl�-^���	?�t6��p*���HA���]5�+ȃ��+���)lV� �*lջߓ`�����s��M%Vy����=�pUK�E��uZ�(�2�A�0����TG�{��ں�0��c;�
��/��7-0��B��=�;���y�/�:�z���^6�HE�g�,+����������Ƶn.#pQ�%�`��)����L�m	���Ri��P�Ϥ�Csa'U�G�2�ApY�5߰v�u�϶a�3���� ��D��ߵ���� ���M0�D���֎x�<�V?�����ea{J��j�j}���h)J�R^G���!6ΘM�
�lA���r�'} � ޣ'�d�'ڇ���`�{.'�N�فb	�G��ޏX"��jۘ���%)*n��WtH���G�?w[N��]eL�KM��)�6XlxVHYEB    7265    1660�ٟ�!�*�6�i��� Mdl�����g����% �ߦkQC��0~��E�Gh�Qj:�OS�\I�u`��7�)x]�n6bAZa=����������c̻݁֕,@�/�.���a+��蜵��*Uˌ"r�%����S�9�k��1i�+zP#^I�2��2�a��qAS���}���ұg��"g3�.���f[H�	�(��?w0<�dv�]B2�iI�Y�1c�����w���9]E�A�`ES�P�T������Ϩ������>��07	�TH�/��[�.	�o�Z�5�[�v�	��'�����m/?9sA�\ٓ#Q���WJү��-�R�'hJW>�$���~��P�Ӡ�y'cN�-[m��;��~�gs��iNO/މ�,�Ӌ����𶡻tG�"ʩ��V<u�8s'�lKpܾ���䐿Oԃ��:�"��d��~x���f2x)9���ţ#�X�U.0��u��B8}�B���XR��u&��7�e�`|��%����WR@��Rm�O%�K�X�_eO��!�O� �dS 7Y�(�jh?�1B�ro&(D	���>≣�c��.���zJ�y+�=u�-�s)�	i��e����_��H�ƅ̷uo�u�!�K	��b���<ʲ�T}C��YU��๓��RK@I?`�jn��;�^{�^NgӤLy	�s�U]^�����]���=2^�,�,m���Tr�����u�W�!�s\��ݚ������Ck 'ס�?Qп�gwr�/�M���/4&+�	Q���U����}�6rd�B=�vK�M��������Gj�7x*h�h�>�e���h%6Ac�}{���M�ndG�=�4��Z� �_���&�[j&�l�V%]O��n&��M+�
��L�+��_ ���{��W�`����HS�l��w~��L�/L-���H��w_�@���Y0[\����[�1��Jϥ��&*��=˳�O�&�����+%ږ�����L������=b_�aO���٪#b�ߜ������q����kf�2�ח���=)䊣�,{�KZ���o[�{���ub���#W������ȚE�)�Xt���z��XE3���_�6k��Lv.���ewG��B+m�%�۸l�pϪS߃"�+��պ�j7��>$,�s\}���KQ�X�(Tg�i�a֗�����3���>�&�=�6�l�L9U{QM�0@ǈ��-}��BB��1
��l���R�r�j��p��O�W͑���K�ДN��:�.��C�lb��I�4O9���K�I1qu�pq}�:�'x1��n�}����6�����aɩ�O�J=�2�]{jI%4�jM��: �0�_�fu��!2�u�`*?z�>�����+�v9)
��+�]�p��E\ssl�K`�k�����߽T1�s����R����f�U���>����W�< -R��w1=�ȽW����/���H��H���0��^��$n��4�$�Af`���>�l�Uw��K>��Q�'�1B��^y�K��b=�GW�wjz,T�*C�#�]m��W9�|��<��r�ż�jN�v�Yr[�_���D�h����J��&�ըa~�R�;�8#�|�sz��cl������H&�PP��|D^W�����f����͜]�Q��!E�#��P��M�Ty��s޵𖻝��j�w�%󐲤�;��N��c�p��s)���Xᓆ������)�H���5&�c�Z^��xu?Bɇ��߬�����e���
{lә�ږ(ٙW�y}c��r$U5.���w���=�)�'�{"����L�Ή�D�e�;�ε#�3�#M��	�����z �����F�=���N��,�G"� �週jB�]l�Cx�5��U~á���+]37��(���h�nE;d&�5��̪�G8������X]�:L�([�!Xi$��m+,���}>���p;�I1�&n�����[<�ʝ�٨6!��w��2�����h%��Nuw�.�/���\�[�B�+�'��;^���:!X�M>)��ь�-�|�$��&���(��R
��'b�"��XV�����%�$��&�l#/L ���v�U8 �p���M�(�8��@�j��(ل��8���[�Y:Z3_:(�ܰ�f2�/W��b�4 7�����Ed�P/5��υ��C�"h/l�]���9+j�jj6�bn�&j˱lt�8��{�gU��)������c�m��?G]a������V��H��%�5�Ӳ(�G��h�J�_ ��<��a��et��$naO_�k�}r��qJ�v���S�V	-N!+����]�5�.�+��E���㿷����^愛B�-��6�d��_g�=pG'H�E���>���
�,Vn���W��9���b�r��0��e�2*,l��E��7��?̇�)����m2(lw��=àSOk��O���V�R��&�xx��Q��x��t�W-��T<-I�N����]H�~ݘ��s��V9+u.K��YZ|�u���P�kk%��~��G��AXV�z(EP��|�j��[�*%ӹ{�������g���$�҇B���q}v�Dk�a�y��m���K,$�`�X�x#���s!�K�o`47���L���2p�=P���`��xIu���u�VUn�QV,e�\̵�D�-���7��RC�v;�eU&�v!����>� �.��"b�1�V�'��d����KP�s�z�̭�o����@s9 ��&>0{Շ��ֶZ� �<}���Ŵi�ej�}����Z�s��g|r�zV_G��ߪ[����e�Oa4젧
{�	�΃Z�	{1��,gT��3�`z�J�5�Ȼ�����3h8+������|�9��P����8��B3�L�s
~r6�����n�ǝv��1�$�/�����J���������l�ۭ�rP4��ƾ� �A���ݦ�C<�?�� �X�D������7W�{��c�b�*�h6y��fҚl�i���Q@��/�홃P�^U�2���I���$-���7�޾�[+��Q�ŉy`�)φ�t����V�m荣�$�4ze<����NWU{6�>ig�N��q��\7r-��#*�;� ������m���Ś��<�o�7�7=��QTIG8��Y9�s ��j����e���I/eR����ߔ�YS&��-��ĉ������t�0��`O�V��.Wu�4V �p�+0�E��J�P�O�hM+��Fxuɡt{M��� r��h����yHqr&��.i�Ӄ��);А���q�
aA�L��'�
\��E�������Lq��e�|�������LT�Ҷ��|�,��紸��ǽ�{�۵���K�|D��+Ad�>�ى�>�����QQI�� �D�!mԷ��� ��a��S�O�\�`'1/�����4���2;P���@�������0�͢M�I|Y��Y/���0��M��>'�Li�t�ƽ�ƁT��<��?н]�-����D�����FuG8��Pb��Hn����q�˧��lZ��x۠a��e��P�E�cl9g�F���M.�}�q�7Bȥ��<`�zDw�f*k�;�B�A6�����L����7��v�S!��� d��.��WU��i�����V�l-����$uѯ������5?g}N��G�6���5L���:����S��%AB�,`-���ٛ-��)$�n�W�
W��`S�Vgp��ER����4�Tɪ`�ps��+#��~O��(�[���̭g�iH��8y��q���n�8�9Fpa�����0~E�*UGr�:�4��b�!�yNR�B4����`��5���#�d�P5e a0�3�x�G_�xi���bn�݄M�	A���/K2/�0�;:�cF+^bL�@W����F-��MK Y�gdA�����<�|�=��U��̅�3cF���}��!Bo$�7��;4-\-N�K ��x�O�R�,�����舟_(�s��j�7�B?�9WR��~��kv�:�&U��.7DD��t(
�oa���㊛WO^�`i��"�Da�f��P�u�����풆����GY"@l�5iB~�	�s;Z�]��'fR:z:��IC��n�IA�:yɍ;�����!$Yxb ����gV��ҁN��U��4i��rP�0�#>U����-�{�u%����}��:��W˲E�����9j������<�Տc���D�hC�.Ơ��<ۧ �C�_C��,�M�xw�\O��=��� ��:o˜�R@�n����KoP����_@�C�W(t{f'e�i��Nt�a���Ω�+wy���A�M
��W�"k�"	����B=�`��
����rJ+;�Ȇ�H^����U6��x���	��.�.�Om��)�2�$�v���������C��gI�%_L�ͤ���=�FG�H�3�BM���B$xâ6��	Dt��NP��ʡB�=\�-�-����BD�lCx���]��à��(���d�|�S+� ͱ !|ez�Z<~v������5��uc���U�;D�Nu�"6-���P�K�W�#Kû����:�0{\��]K��wձ������,��{���m�wQ�D�^�?cjG�Y��y��%���)�^̹glF�4҈�fܞ�2mx�n>[A��g{�R~�)��k+��B�s4j��iZ둻�����V3��߼C�|��2�SHh��bK)L��`��,=����%sM�Ho-C�d�m�n�{�%b���|&�[f`Ȧ�')ts������U�1NĊ81��;9�@c�Bx]�����B����(Q׌�qFI�kS+�).��r�D���B9{�u��ܰ����Ͱ��i�S���$e�(�̖A�O��q,���+8�bf3 C�E���¾/�d�+ː(�,Q���}'z|Ygj:oA��I`�U����pGVB����p Ԟ�R���y�l�Q�G"�)k/+�u,>��Ң��x}�w��Ӽ]4���^}�-�{��8���bL릡8pB�1*�w�rl��w(�8�+Ef3��$���"?�J3)��7K?Z�j�c׮ꝭ���^F�e��	�ZXGL�͆�ہ���w��)�K>���_:�y�-:0�����{���
Ǻ)��X�2 ���5H��k$G1�LA��X�56\VgΌ,��!�<��ȱ*4h������o\�|�k��D;a�A#D\$M2����>�`����Z���^CM�w�����+�96�_���Rձ�����3�	�s����~����M���Jo}8�b�@�:�AP���ٱմC޻�_��F�R0<�)[�S$�+m�qs����
9I������x.��t܀��AE`����d��H}���{:�s�*KR��L`�|�V)�ٻ��#"���G�^[�>)���A΍�C���.��E�@	�W3��$o�7�I��B,�BBy�#�#���4k~ϝy��Qj�WS*�x���F����0Ō� В�M��\�H!ל��E�ϿB@D���s�1�����К�E9���C�K��CW�wYO�l�ܶ8�U;.d���i�)���Ȟc.��G��Wk�L\f�P�H��Bs�1G���[�ª�B�.�4	�M-�Qou�H��r5�