XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��)�$���z���6�;�$x��d�0�!�k���m?r�B�Ju�^�P����#�OO��2-��<C��i#�?'��,��?w�7 ���f�x�Ӌ�b/�M�WCp|zҞ�ū��h�;�
*J��ۨ7��k󑂱�-N�17�v�}#����)k<�ܤ4�I���i�R<*�
j3��Q֬�E8�!g�D����H�I� ��@���@��=�b��=��	�e4iR���A	a�Y�j�.@=�?L�q&R���o �?0�j�j�wI�<O��F�A��V��X�\����V�X8*~oQ<� �('������p$���'M�������$���)�	1�=���é��ك�su^�)8q2L�xX�n��\ͼmtni�χ���`�'�iy�xr���m��v!�	;��p&���QȰ:�v������7#�$7]�T�M���R�l(�xa��Â������J�c���;Q�����0���<[gs�]tS#lbQ�_�9�VK�t�4u+�y�"@"t)�q*SwT�� A'�q�q����j��X"�"�~q�Jݓ��u���2C�ɐH��Q���e�"�w�����A��<�'n-t2p�^��Z�f�����.���G��C�Mv�}`L�������<⣀�)����ۦFJǲ�����[�38�1��\�*p�J�KQ�{�%��g(���W��.͠��3±\(\��_��d*p6��9?�g8[-�,�'���XlxVHYEB    9fc7    1fd0(5&`3+K:]I�/svI��;	1���8��ʴ��TR9��<HPO�]Z��Y�	��SP�'	hMQ�b�^Ӱ,=[��M�o�Z|�1]eԍpU262�T0�`��v��\�q��d'��ޏ~a�n��N7k|>�����W�.�s7�}��q�a4e���p�g�#<P9L��pp�~�9C{�>���{��i��Dq��bB��0��R��nd�>R6�p����v0�-�U��|l����p�=�Y��X(�kZ��hDjT��/��)E��H@Z�$��h���iɫ�yI�G/@d93[i�ib�7�΅K��8���Dc#΢���&)OqJ�Eע��� \�:�`���,�<Ǵ��)~��\I�*�j�q�e��Lm�n�İ
�W�(����ݥ���U!��;��}.�S��MՁ�|<�21���.4����O"�4l3��je$͍��"E�F8�H�١�>���j�����+MGL��N�a�J�oԫ�L��jX�xx��]�P�;�i�R�TW�u�6�O���/�s���OXX^�$ (��Y���Jc���}���Y+I@�D��ΦQ䖑�$���a�b�/����)�N�\pv�V�b%��MAn�Ly����νG��6�B��E$��׏��~f4�ΝD<c��\�����©����u�Eޖ���EΤ-Q��R1%��T�����������=fG.Fo��eu�Ւ�@mr��;꙲��yXj�4Z�te��9J�K9��}ԑk�a)b�*= 8�Y�j쑊�8/��.�4_ݥɺ(J'�Y�swz�dB�0wqt�j�����~H�a+H��݈��j�R�g�x�]���+ɐ|�}��خĐ�t�
w[u{�E8������#,���K�!}�~ �����7y�P��oTK���s���8�~��5v�E
�����}����X>z9s��_�Hߐ�nq"0��oC+|U��#�j���gb�����@e��<�t���.�N2~�6% 6߶�_�&L����>|��C�h�h�7�����wJ��Arv�ʉ
�wV��]�`��b���������+s-�#�}k�-�-�����k����ƌ*E��������Ħ00��
��3�q2��}�iłLg*ؐ��r!���uۀɥ�5����:�����+L�>3M���oB�@��{eNP��I?%@y���O"�?�(^k���BLs����h��oO����}���l�m��~z��2k�<P�[d�1���х
Dwc�ŚK�~�u�� Bd�3z�&��p~j8�U=����p3O�Xp��V�g���ڲ��%��+;���r.�m1-��e*�ɛ�qzQ>4�T��[�7��P��i�y5{�X��7��k#��,������W��);y�
B?sM&�� ���a�#�ǜ�~���$�l��SQкѝ��k0���m5�{�<�Π���2j��������&����Jt����O�r��䗄��e�����k
�����v&��΄c�쮏�.:�r�L�0.܉h�;l�r7�FN&�+3��)�uP�QL��tkK�0'��ẹ,��g��5�1?���kRl����)l�k�z� ��`�FG��⾃���mݤ��Z��|Y|&D�E�i@�/s�[
�7k\7Ē����X�����������Q�o��\�f��YW�4,4L#�
���{YPS!�ԪK�zl��Z�Jʻy���b�꾡R�h3f �[Ԟ�qq�afn��0�f�~��z�w��BG�Etx����he�2!�ƹ.f��MJΜ���跳*����暡tB��p6�:(��f|�<�D�J�����4�Nm���Ȍ�!�i��ᦗ�JŪxP֥J����{Xr,��>=K��(�'L��;���w��Vp���K��D:ܠ�y�*`.@o������ۗ���V5g�](��N�_�B1E�T���j� 5��J�W�c�i�߃��ιlB:��^�eayl�{�ײӦ�>a��* ��c�"�{@y+�t��ia;bqI�%�C��i=�%��A��D�
r�Mߢ����R/�c��>&��MJI~���S"~��%�,�ɊSt�N%�����h:���=U��}ȴ?���fģ�52�Vx�'�O<����K:/l�?ګ5^������~�z����n�@f��p��~>;yW*�� G�葷U�/;�*���)&���!�5����U=�>F�6�;��EW��H/��8����2e̡a�Req�9��_��,���ŭ�Hl2L!l�^���iӣO��2����zV�Z����z�}�L�!�G:��C#���Z�A��ꮃ�i�M�Y�v`�:P��˳��-���2���GR�~ګ�t�xe�0Y5�V�:���n1祰Y>F�c��+���sZ��T�WA���B�G�G������������ v�6,��X��zP��"6��g�F�A�u�g�eu���	[	[�	������IǘÁQ�ZEuę��G�HZ?��{ 
b��>�O_&z�M��4^�B�G��)�>L����R������;r�w/�>?~Y�?x��Z�w^�粀��)�)&�&2�hd��ۊ��-l�ez^0Q8�&�,_�|�V�1��E<��w���v�Wχ�@��.��v����6�=D���tw�h��I��{���O������0���R-�\���V:�i*6�=�iN�����g���v!�d��aA���!\�����-�Vk`A�hnp̏��0�}Q�k80(?I�Û�ϫO�f}��h��w;�����#t\���@���gf�}��I7��2Iu����m�Ɉ�:��Ȇ��9�@�e�N��q�O�R�����Yj0+s(+��"k`?�a�aB�TAG\�v-OM�Y鄷߽5��,:pU�����W) ���D������	+�e���<pFDN��c�G4Ow��D�E8@��ܙ�	͉0"��D���Wg�����yI�b��9��d�<&]�H�Ԧ���X�yx��vF���ny�-2�r��pa� �,��.����נ�;� �@�^ g��f��A�	��	b	�a��N&���	�lzM%@��n�QQM�Q�Er�H(���jJ�������Y�=A��6�_g3w�[�,�>qе<�l|�Kp9�f�Am�s��EG���Lf�9�ά����E?�,��"����>8�^�N<�sx#E�	{�g�8����k�����OZ0Rvc��&h	�A$}F���j=��=-���#m������HW��nƎ$�n�)3�6C)PӺ���r2{�}�;_�������ɻ�}�28�H�`�H�$F,�&��d\̒��_l>��&������A�|7q*���Èd��$"��	Ӳ�G/���.��=��W�G�&�=��dY��S��ۘ��}��c��f����=p�������=�D,��x٠ޯc��1�0��R��K����3y��/��>�$@&�9���wV��K��OӞ�p������ݭ�:�!�v���ؐ�vmgv��_I���z��JF�1����"\������ERL�+�ׅ�?8�t����JPu���O��Ғ�;����<t�\$:1���&?�!+�򵀶�Sm�J����C�-3RGM�_l�� Y~u��5���� �P��!+�y(l?���"�2�@n�)�Q��%�ee�b5��eP4y��3}����Iց�h[�4/�[�������Ώ�ʥ�a��;�,���\m�BE��ʁ�XW ���f��R;�����q���p{n�)N����7Q��(��j�p&%�x��
�OP�ʆ	SP$�B1�U73yZ�|l�aTv�J6ݬE�U$>�W/��к=�*B
�|�i!O�K��0U�IIR*�z�i$��Ba���e1�Pm=e�/��jҳ�d�����[}�k� /�i�ѝ��)�-� J��vr{�\2|;��׿��>��?�ݼWM.5��R����`�?��i�����!�T�@H���o�,V�=+p���}ѢO���5��G���e���������m{X�:S�������}Q0���z��F�� �s��&En�X4~L2i��D���x�;1��L�
�g����O?�=F�0<�#+ɱ���Z��0���#=�&�Vj/�]8��S�`8~��O��9p����H�Lv����o���[�忧��(�������`s�5�V�s�w�o@���Ļ��+|����o�h;��!KK���2!oĸ14֛����bi���7���gqh���^�K`��7��f�;B�o��H�?��f�����f��6o] �0��A�6�%��_B�"���k
��a
�V����<�Wν����3��\{�A����>���U��}�����}q����<-�DL�Z ꔹ�R����Z��! er_�g8�HGQ3bF�rY�,�a�^Tm#
T����ͷ�@��mO�|F��8_Sɲ��6����g��8�����%
���!$7x�l\8��P�\'w���WeTw��A����ҡ�J�%x"w��v:��\�WV�9����|�{���Yq�.UA[��ߗ�]4r���*�DLE�B�|WA�þ71T~�X�
�*�P�$�F��p1'V��Dg:�^\]��z���ߍ�.�� �+���A|�����r���zwu�#p�

=xn��'i�+n)��_GT�[#!�^��B
xa��{�\����
qu.�Կ�rR�ӼF����#$4�F#ǡb�h�v�����>��5s�z�{-�F$O~�����,�����'����H�f��Ǔ��N��uB��5
�1 �q�n���cCŧ�w��}�X��t1H�5���&^����m�
)�(Q"�� ��JQY��y&����-ê:�R!�J����W���P�.�w�$I�k�N���u{��}�ԧ���Wv��X��7�b?IK$lPi�� ����H�Evfg4�y���l�����	��<���:8�Ŷ�&����Ǯ�������;{�!n@���i�(8�z�U�,�f�O$���i-x�F�A���)�|��H��R��'l^�'��}�� B���@l�&����>O�d(BY�Ǳ�&������aTO�i������<̎z�G@A��F���%�Y�����)({����"�2w5^�5�?V�E�އ{u�qcL�#�\^v�o�,ZQtW��ؙYp��%h�_���x�?�D�w'%���	
���l�.�A`����� 7dץ�J/�,���p� ��?=?W.�8	�?W�������Z��2٘�
e�k����2e�9�<����]G���C���\5�	��.�D�s��������ǅu��M�y�y�t�=�۝���.�L�s�|X%� �D��/[�E���a�7 ��r�ˉ<	rk��V���1.ZO�����k�J���F�'$�7�\\�l!-��2}f�"C�#Z�p��ơ�J�ȅD�묊�,�a�7[�1�Pnu}�kb>io�ӄ#�:���]̄���=�G�9�i����҉�	_�Hþ��q0��|L���t�z�QM�c�@�]"�X��灛�ҭ��[���ݬ�}�[*�mw� �����(Ġ�u4$���!���= ����MA��KX0���@�(�������a�>:냩���[WT���%���zr��QT|"8�o_��"A�P\�ŏ
:�j��Gx��x���Y��$׫bx0a�a�(��$-w`������pek�J6���=�L���o,��lbJs��^��Y�|(&H���]��A���@L�uM��C�ӓ�S�#�C���+�[�E�	�G5�ux�EWU��xXv�£hH-@��ҟ�ۖL}�a tb({���}��7zv{4
�H�1�-GpX�L� ����x7�4�K�@iҹ-|QY78� {S�1�E:N7��R��4�8ʮQ���� N�E��3v=7���F��}*;ū��:��f�G-��_	E���l*��Č�+���3�N��(p|�p�y��^���x�I;��Ղ��&��c�=�#-�n���M�T	EYrh��u�L4��	�6?�2o{eaW��A��Jf�@�+����>���C �uMD��
����qV��+SP���w��u�g�Ӻ)��4s�ywS��f��$���a�I���3=c�R�w������4t5��x�#
�h��p�VCs�شFS��&�|{�c��b�4潽�@�L�#P��z8
�p╦��>A;9G
�h�s�(����(��l0�\~�y�S��'SNOj'�w�EADm2h\{���ވ��C|�H���D劌��J�v5���~�R�׾ٯz�������c�.An�e��MM��Gϭ=���0��A�R��u��x0���ƭ��.|�t���}��uW��.J��Ք��5{m!�y�ਏ� krK;R��(�q�ٯ���gi>n�O#��/�&�{��f���U��� h~�k#�ԩ����\r�&�l��a{��y��C��"o�#�r�,m�BN�.�N�E䲲a���{��M�\�Q��n����*��_"�]c�2+��ӱ�����FX�Dɺ�;�w���/f)���
����g���g!n�\(Ǖ�(VC9� 4n�!���2��������6K0�����m��q�jcx{�h��6�À�
xja ����rU3�����X\�:<L�A)��,�������P��dp`4�ۿ�^&9�+�A���[���8@�j����2�|[���)�V��g����J�E�u@^4
��ad2HFAT�Q�W�����/_9�d�]:�W^iC��d�m�BM��2�qX_UU��9x���S�vx�S��j3�&p��%�/�ȟ�l^�Hb�K_��%�����^Ԥ��Orȥ���˼VnJ[ ֮�k{yQ��� �� i��MC�RL��bDʃ<J�nq��,�ĝ���5B�Ӿ_�6-��~",�e�)#޹�xA�9K��B9�"H��^�J�Q��3� ���i@�`�d��bs�%�g�8+�W��?�h lP��ltC�t���J\�O�3�^�)�?O�fJb�\۱�h����(_���%�yS�SYw���~�=~N��(��������� 
U�P9�Ŵ���+�=ei���^��	�t7ک��g��2|���8��)���%R
�^��K�(�	��-K1fB^�\F���}h0�2���ؐ�/K��2#ʞCV�#�dH	%����U�n]t9��f�'h��x(���'79;[hO>q	W����-���R���
����.埆�=֩�u]�",,�+ǐ�|}hJwë&�`T��Ћ��"zT�vk.�i����,���>�z	bQ��<\�U� �Wܺi4sj�"J	�&X��>���d�1�@�(y�x�`[tU�@��P�vth�'a�E��<�g�͊4Iv說�m��h��)��b|����{�W�ڴ[�wR���Y�}z[.���zm�~wD0���C���s��_;F=�����
�:8u"�|�c빷���.�r�{b����0��� �"�⩭�3���qEʧ�bd�Bc63���%����Ϫ��0��Ino�P�
F� b����4�5�Y������ ���a�b�Vl���\���Z;�9��Og~G�~���'t�M}�����y>}Ү����뮃�`�y�R֨���春Ew����r�b��v�̡�8��#%E@=����i�bH�ѫ�c���Wq
�i&��R�k "��A�8Jv�������>�t�_LEC1����
��1��8-�p):����^�W�[����UM5H�(!����	k�y�*����!c-�jVB�Zue�dk-��y+�V�h
�=d�ڸ-H���D�]Ln��l*�Ya���Sr��HB�� Uo�dEқ�%j��i��Dv����t�?e��۱��,q=�c<����2�8�
(�TX���0�`t��=ۃ�v�����Q}�F
E����.m���r&8�