XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��!YH������ W�7#�����}�mڎ�����k�X�U/���V{j�
$5ڋ�^�.��!r�`W�4�շ� �Ob<N�A��+���/��-ܔ#��@Y��=�
\x�!�.OA �q�M��x4Z�76��?�UW�z��������9=ؑ�=V���U��B�KPP`�U��g�FI�$���Wb��v��Н��;�gj��s�:ݾ�IuPNbu$�1m�_��_t�+-�,>b�*��q���4�X���{䋱\
�X_+�[$�K�qY�b�����_�01�^�������s�N@�>�_Ǝ�ܺMq*4v?<A[�,����lZ�|o���S��d��9�@�O�L�|n�ڟ�}>�x��j�~��Vdx�e�FZ�j)��S����C�]ƓXèo-,V�ohN�u7d�e��P�#`�/U~��^`��B ��6�f6m%�Y���q�,�Ö<3��&\./�~��T��v��_"�]����Q���+��k1��I�$��ޞ����\�e�mT�KQ��/��L��ڥU��|O���33
!�
h�s�i������\�(�3�Rh�$L��1��R�k��*;�fP]���=��$���?���Qh����]���z4Tn�	(yE�G�}6V"����U�?��[^Q���Aw���s�%I�+/��P�M-c���\Gn�s�?���pV���� M(pbnR�E�S�@�;^ýP�y��ہ�>��XlxVHYEB    5224    1740�=���1N���rҫ�{-(��	�^������+T�S�G��\�m.�\�ǁB.�������}��i=Q����&�W����!���Zlj\	{m��1�\s�9����\bnqN{JZlzuэ/��EIsh0�mt2�Q.�'�E���Y��^X��=��.M&Q���A	���d5���I� ��G���y��I�{�����}m�\(�0��Z��!3|5]� #����8/I��eCZG�F|�mC_$�=ϝ�dn�I���i*�q�;���%>ăYן��l�ٶ�D{�O1�@P����,؊3��@�jm+{V�/&��;c�4��/Z��]g����z�[�c�7��qՋ����2
l�l8= �U�ͣ���g���wD_,��f�����i����������W<�Z�|�V��g)3˦!�:]��&g������� �l������#�Q�ԽD��x�"m��}��?��r�V �i�*�m$g���'io��L�AВ���Ә����DJP*��IB���`ᆆ[�,G�JV� ��$Px���]�Й�]�� 1�k��U�~��ƥ�Z�U�]�Q��H��J14J��I���)1X����?vJ������k���"[�t���rsn��qm�8��0x�w4�(=VN'�5�f�?�d����0B }/�aR�~�6J��}tY� m�Y�kU��������M��A<�G�y&�СҨ�/�w0%�P�ݫn��4y��f}O9}*WF�8����~�g�*]�������di�����zv±����3ݍ�$Vƌ����
���>�SR��b�
xt�`��d�g����1�K��Y�/{\��v�vE���	���3���p�����TR
���&QB�u$��ӓ����	� �������7�{^�1��P�cr�G[V��?[��3x� 	�0�jN	J���Ϩ;���IJ8}A�a�L��U*�)��)��SS�(�A�6�[d`���\���6O�=�Q����6t	�<@#Lj�����VoO6#�p��	��a�}\��$DW�2�L��p��iE��S��cG�0G����W:c��k4
���Tv29�)�[��	����D�"-��G�>1�+*ک7�t��f%r�%:��F��S�,�G�afg�A;XFs���%�t��-f����;�]������0Nf�E�j���&��~��$��� �f'v8��8��7��������e9y����^���_��� �����4a��v (�#�vl&��i�=���(0� �?�Y�E��78&��6"��	�^.�F��K��l�f�`5q�+-{��&��т��[��ŝv�,��C?�?����'sǳi�J�7L��HZ� ��*{77���1z����K\�l4���%�G����]�T�U�������9�`^L��;G��|��Y���F�%"Еb��ȩ���"m��h����l�&LNwI"aUul!���5�Њ3��r@��ᓇ�Qi4���0vv����(����;ϯ��{�Վ4� ����+�N=�,���TGAғ���c��+Zа{3��=D��y5�j����� 1���:���Og�:�f���23��i9��y����-������8�8�Hr��N�ya}pɻPhG�Ars��ؓVf�A�!oM���*�<�ÆM�*	�XM�y1�;'@H�.����dw��+DN���C�	�i�`�R�Gߨ�����#/�uD����5�ot�1t8ӥM�x�R%U�&�lR9��ь�S�O�ڟ������tE�B��(#�d7��@��M���㷗cb���� �RwgcsJ_f�D1 ��[�"�T_v-�!P3=!�N	3�+r��ht�����36B�e��i5�h s衅e.tË���y���2aj'�$F���FzS�Pt�Q��P0����G�}oR���-�k�h����&���X����4��pZb���̐t�-�ܹ�J3b|�����2�څc�s��R;�/?k�4]� n9WoI�	����'75L�qh���d菇xyؗf�V�f��e�ǽ
�Y>�JpY�T �UO����5A/����[�}1
X��a���P��/@��� Bދ�	T^�.�ւ�#�}��ZS�~�c=Aˡwا���(���k�L�fA�����p���t��i'�C�(�q��!��@�k��sR�����9���F����,I	q�9�5��8<O���6���i�{���ʩQۈ>�*K�X��!
Ԃ��+��ֲ40Z��*�T({];�H�=i&E�D�ͤU2��dW���t�}}�f��[�h�7�����|,\q��I����󶫏Z��e�i��O+�Dq���߭�ߗp��E�׀��R���K�#��j8~+Uc�� �uG�}��JmI%l=/l�9$�����@g�NW�H����*DD>��x��&>�����,�q=w���*4~bN^	�
�^�W?(����x���; I�Ѣʢ!�����p�Pug����78�>L�����T�F-12��<�f�CE��n1LJ����i��"�ԺD��T$�`���d	!�e�1���9��e�@�'+�pM`���k	���19�Q�����)�ŏy"ee$�HH����_�l���T��!�U^���%v�_���v�KI->�Sa�8�.:��ڐ`4�����Rc�/S �;�X����@��w��m`-h�N��_���9����x��t�hQk_�q��ڤ��A��Q
�B�+>1�dNG9���6�g������,�z/`�p�,�h/��u-	B���r>�}���.Ӝ�9��$��qA"�����k#>Z*��,�6,��t�xIvi����y�f���Q�5
 �����Eʧ��*�9��� Ų�~�O*�2!Ѧ�[^c<f�L/��@�ICA�W��Ϡc�DG|-�7�a�ΰ�~���M�e��������� K����E���J:x�'��)��L#����lL-$e�tk#�e�<�_�K���\����l���
}=W���e�/�A�m3�8:!���
�����՛e�Y�b�$	{���^�0=�txY.~�٘VО�176�\�c#Z�
t�e2%��*�!#��D��.In��r"�P`Z�i�3�bcqchg2��)/q��aII���& �Ɵ{�2k�3`=w�#�=�A�\�m��}R�@�8��rȦ��Rɼ�R���l�S��ġ���pD� ω-�d�'�s�s�s�3���*����YƦ,G��=�CA�Z��`@����p4��r��y��e!s=ћ_x*J�cfa���s��'x�pѯ�4w"�	�rt��鲤5�5r=�,l�u���ʖ���T�UC�oO!�~NH@��m�G,iJEy��gD�f*���pԆo���Mp$XQ�!�2��f���n�}?D(��;	��wB�͆*"�ч'�I����L#�p�_�m������38���)6#�x��E�d�?�d�``��ul� &��cepV�C���(��������=xīDz���Ȉ���@�c��R0���_�8N�5�0=�9�1�@�+:��� �b1MP��$�!��^���j�!C}�dP���C+Nd@�^.[���J5��p[N��!��0�I�H��h���a�}��
�>����f��5"��z#56X���#Cb��D�4��σr�%��0ׂ@���:�����{iO.�k����b�|��}G����+��2/�Nvr�_
�T�/�M}�c� �b��x�D;'W@�|�0RE�2�{FV��x^~+�
�g�M�Bu�P�F֯ѬοBMG�0�{ȝ	�?�j�-9.��g��o���Kf���o|j��w��	Hh�a��ٝ�=���g���n)s�E�8E�씻�)��~��x��4A�8�R�*^9hgn����N)T~KvJ�e�׾�b�FF�iSt7PD��E����!d� ��`v>;=Pr��~}{�^�X�95n��&������V�5��6�����zt��{6N��*x鰀���		�m0f�d�l���	��dP�D.ȵ�vS��O��9V[:I��]���y�����|�%J3=y�)���8,���-�t���S����\P�(�i'�a5��C٘,�܋!��_R�ޒ���g25,��*!,� �~~F���5�}�s0�,��(��3G+��I���9���U��d15�e����a�_�p!�!5��),�_����(�y�Y�	�\oU�I&�.���E�U�J����K;�VS�ԉ���5���8ԫ�Q[���4�ɸ����	j~߉��d�R*��FZ�G�@=%���u ��z ����~]����$�E$����놄A�j��{���.����]�VV�� �j�~כ��ƴmvU�T���2��|����$"o9�"=o~��汻��w��@P~@�n��IAK~�h��+�zS���^`�KI
f��mb��JԨ���U(�~5��^�J�{,�l�w���H��h��p�nCY�2�����e5#"Հ�n�z�a�,�˵&������l����N����;�t�����ED�������/Riv-��-; �p?�u�ڪ��	�u�	`��*��wZ�����-�];�|�n�ܛ�τn�����eR�$�f�m� .���j�iرSE�Dbg;w�݅�Y�6푳��g�lS��nٖ̟��^�K�����B/�}(�����x��,:eB�$�&�@�5��b}T�8^�-�bǝ���Pt�S]�Ƈ۫Ę����E����+ptk�����d��?%<_J[*'�T J��y�P�E�u��a�;)ύm5��o,T��<�H��@�O��sC��iA�����1W�Zh���H��'���#��Y�cu���v���3�<�<~�d�
�("�-fK�x�Ri'+���T&�$��t��S�[���M�`.�ie���8�L�{�c�!^��Ο͌�k���T�����tfb�ab6� 
��.\bƤz|�Y�l���;=0cހ�'�&#��.�~��s
�}�6�	v�>4���Mk����^MM���5��ۑ#9�˜Z����/��թ��נ�!�P���d-�})��?� 0O��>���@�4��q�p/�8+���_�bD��_˂<dկ�8���P$��ά�8;C��3�Yg�z'f"Uۿ6"ˎ��g�Vb���4��Y���/�Fu�Z��AD�?Ѭ@eT�q�y��ίT�j��Q3P!�l+c?��:J7�\*n�$����Y��Ʋv�'\Դ\�6��z����d�F-�>����6F�N�����\�A���]c耍þ��z�$�<f���.|�@Q��^>,��� �m��xH�������t�f<r�9g�;�B1������OHDU��Gdk�	�x���� ���cu&�Ժ�K}�@堭�1�3��u�������UG L�u��k9��'���X����R��F	�� �{S\Ɓ[
��Ơ��N�|�M��*mq�U��75D@�kEA6z���� pUs.4l�̣U3����#���-$ qU:"ru)����hB�6EP������ؿ�6��S��t�a��:�>��Wp�:�q8�Q���������B���`���S�����Fcݒ�X�ڂƿyx�Ҳh���'ςD���G�P�ѱ5Iq9��������@�������:ٔ(h�>"�jѬ���Q���+i%��C�&Gsm�&o��c�}������mQv>��N ���c���Q