XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�������0��&�9J�R�c:l���̓z��X�ل��,a��w-1^x�����Q����}��&1�ς��^H�^�Ǔ�GɋĐ-��q�h���FW�h0��V�(�'��6E;�ƫ��+���e��&�j�������z9Zd�����ܣ�1�1�Q�|r{"�w�����2w����R��G\Jw>�����CjWRS9�}w)�]ح��$	fy.dH�u	{'I�GM���i`������~�q�ٗ�b����&�0ڪjz9]�k���
w������?a���$)>Dzl$�S�7��u��)A�� !J#�O�5���Pgt�V ch��%FT̭Rw�gZe�;����D `B�հy��c��.��?�I���M���!}*-�Y�W�[1�_⾥�w��= c	�
Yg&���0�	����0Ƙ|.�N�O�%�����զ��S:ܔnr�F�y�
��$�,��=����S�aJ#Cnd��b͟��T��`��f��n�5�+���}�6v��w��ڰ�<ud6�{W�C�B��1n���h��֌�.-�#�.Z	CT��-�]�a��7���b��2��鶂T[�2UU��'����+����}�ڛ�r\��b��%NX�p��h^uu]{^CR|�;3��� ��w@W7g�'�p&�Q�O��6^�V���3�#�ċyp,�68�g<�W�0���Q� <�O!.���`�#H0�	X���/�t��qɌ1���PGJm����:,�XlxVHYEB    fa00    2040��N�E�f��q�jOJOR�Y�]���":G���M��&	�s�$?P6�[�K�.��ĆQ^RG�3*��-Z�g�������o��\ p��m��L!�ź��Ue��ca�����/;v4�\a�Z� E�#��V���ܤ����%~�&�=������)4?�Q�`� �Ajh��9Ls�]]�h"ẖ�!��q��=lɹ��d�5��r����kY =j)���u��0����H���������w�묑=yz�|8)*1��9R s���Ԝ��["&>"V��V����|��V�<:�+^K����`��aaSxer$>��j�٠۪�[�`��fY���yp�*Nm��`�W�Q@�X�gq�m�~��hN��zňϞŪ��~��ގ��+j�%YY����J�T���vUg�o��O�s9�i&����@5b>a�*4����� -��tY�Ȋ�;b�u�iu️�m��U-, ��V<z)��S�ʁ!f��<AA���n�; �R_"a��j���1!���N���K���V�]�{ ��|��(���l&�Q&��|�,yu����S0��M �R�N�5#��"+��Yv����wu�%&s>F�πn�
o=�\8��j4���_�ߵ�!��sXƚ��Z6�Za�<��_CK�N�_�����*)C� �J����ϒ )��|�k+5I����+G
AdA3�@׼����LM�ܮOH��^�$���6�
�)�-�\5��নAo;Y�N��y!%�A��ڍ�2�Fel^��|<_Hr�j��D�n��[]�H/���OC��Hݠa~A�j�99�eMy��L�)�<���;�r?��C%�ʏ���`��P=.1�(_�&�^��3����>"Ip�a��f=����~](�&�\U�Ö�p�� �:���L{il��B�R(~H�����G��1�C>|�to� �賁�aH��	�R���;��zg(,K�$ܻap5��"]E
 �D&�	��d�������/�A�W&Y#T>Ų�Cy/C��e����DHx��Z��dW����֟�%��K9��fz4y"m��d�G��Q�+���q�
��vS�g޽�Ӧ�	�Jk�&r�9��V��P2�aKc&����L�
kO���
[|M�_+�L=R�J���K��o�O@�I�6_gE�}�(8O;Ⲅ#���=9�oH���C�Fŋ�rȪw��>;;���� D�K��Zߐ_V&r*�3N���ԗ��WDwUʊ�w�9h��yS=d�'o�|�7���>m=GJ.HȘ)�i@,OF�7_�G���h����S�a��7Q)���4�8���Mdu9ע )��?W� �e�:��]��
鿦߹K���ȁ�d�a���s@�2�78��n ��0r��E�,X��p��,[2zg�,!$F��65�o�әOj���"�U�~w�q�G��@����ٔ9���|��.y������ynN�Lrb�����1��5�l\���#m��S������+��k�>���9,�9�N|S[s��y[����g��W*� -	0�hC͒� feG�����	�u���9�'p��mɋ�
���*�=���ũ�>�"�?�~�FaE�΄�LŚ�a��(7	��c��xZ^s\$��B&�̐G���,;�P�-#=�N@7iA�CϨ��o�HU;�H[(��4�e7�nE
j&i�bc� �#w���F{��CɬK0��&��=Ǥ��=��P���@�{�z��&S�Oىx��E33�,�y�4�$��P��P���9Kr3�1�$��e� ���(���|:���}��5
hI��r������5���`�^OU��3�4u)���<� ��K/u��̲�`�D ���b5$0Fd��!r9�h2y�����$�X"�-�����|X@�R��}j�k/e|�s4�قԑ,Oᒔt!N3�����[沋��H�=h,'	 y�*�j"��Ɇ�s���S�	�e�2���^͊���b��y�-3%�׽��<io����
4{x���g�g#���Ge�q�2��~�7[�O�X��MyJ �I�V$(ܴ�<��vf�;\@��75P_IR�?��zU�L�����p��ty�ۉQ2Ұ�2�آ�཰��p�Í�{>�=����t�se��s�v ��:~)�w��J5���VFw��sJh�T(.�Z}��Y�Θ�`9l�}k��KxY��ePK2c�j�.+�C�͎�0�Њ�}R%��κ�@C�����E�,����f��4��M\MՒ,�$FjS�$���@��t���.%��TG n�����p��w�ׁ��V!���$�r��K���y� �tD~-x Z�����i	��Y"�4y��D����c���ޡ�^		Q~��/iͰ!��X`ה��|̦0E%3�i��ß���ڗ���T�(�ƚ�J�h����d+i=��m4�j^�L��"�/����N|\��� ��+��$)"�!�k�MVix+oz�SK�ܥ�b�&Zu?:1;$�tr�!w/���(X��c񽹅�h�|��[���
(��#Q������,	}Rv�]�3R=�7Ɂ��O-3�U��
��3�.�����k
ٺB
�0�`�x ��|��!#�J���i6 ���#D8v39H�u�z�UN�"���`������J����h�K������*�r�U�сF��B �5�A0G��-"��S2)_���2���K	|6iڔ��)�:�%���_R�����M�qWۛ�V�@fS�T����Y�r�a���&����u�(5�"j�ŻJ�2v�B����YO�N}��0�BQ�~��>��?dg�`$�vq�aF�S��]�%"��^�!�6A�Sۢ5)(F���]f,x��D�<CgN�0T���s�")�%��4n���p֖?���Hր�r�yG��/5�R+DCݏ{t+!��O�XJ��9�\��,"-Vi�ɥ�^ڞ��zI4N� 7�ƪLgD}��V�IЏ���eY�!P�q �q�|�����Ȫ� �͵�wOɝ�/���I�RD4�tɊ0ٜ���q�Ýz6��
0'C=$�K���c�A�(���"0�����O�� 0ǟ��CF� �[���tK�4sհ{K���b��Ip�v����P,G�dg���Y4�*t�^?��_�7j�e[VA`��3�d�P��T��AJM	-Qv�����'p�G��c��a����r��k��Xy/a6@��+7�B�ML�_��}7 c{O}���Y��q���T.E:�ʑPL�ٜ̉%����/�t�Z<0��z�I5(��"�e:�<}��KYK�g��~��UD�X:|�� e;em5n}��w�������{�]�#t|���&)\U�
�)j\�?��CG��)g<�˵�)|}��,��	���/kO�k�ν��e�IsS��6�6��_�,�bM?��跶���SD?���ǋ�`1�i@�]�4G���y�:}7&a?7CP���h��4KTp6��`�ҭr��C�������_�A�v��;���bs��+G\�qK��yq���s�CI*9�j��"3|���o�!<�
�pn�3��6�s�����hX�O��r{���j��s�F3u��������	|C�7�Y��K{�c��%��(�6� �w������9sJ�
�_9����uw��0�(<�轵��9f��l���O,�����B2���U�g�&���0�J罉�|���u�&��LKe�$ϕ�v[Q�c��m��St ��/��:i��[׃�����24Oj��c����2?N��TI<1��l�;��E`��?�i]krW�N�o��
���j �0����)e�UrWR��D�	�;U]f;��n�-bK���1,Gw�
��X5��|�#�ky2LL����<v�ef/ה�vT"_�/:�J=&E��b)���>
&پj��üQiQ 
ҥ($�ea���ɩ��j����
U�,p������Ǯ|�\��)_����	6%��;@��%\0�|�L�͊�a�-��e�S&	Q���3��J�/�`3ko��
��Wl�-���/uX��j��z���q��꬀]�U�?���q@9p�G�r�u��
*z�#��L@�����!�l�T�*m����uV}d��i��>O��=:��qǂ���
��RHk��9^��b��
]v��f�"�͹$���u�%z�/ˢ.*/�Av�ǧ�f�a���G������8\��(�Cz��q�r�/�oOZW��O���2�%'�r9� t�Z���#�<�r�MT�&�@��k��|�G`\s��<����<���X�:�����9t���%)��P+�T��	��w	�?k�T���]I�������u�C����{�x\�1����Zo��g? h�<Vb�!�#{�u��r��un3�=ӄ�*�m<j�N�`��k��ģ%0���eM�H����a���|KM�ȯ
jW�)��%�X��d�j�����
����me����Bl�>��TÊQ08e|�"X	�[xE�/�0�3	�u���q��K5x�|��e�cF5}X�n�h) ��{��o���`Y��\Q�����v=F{����A�N�0R��7�b^TtSe���L+K���q �U�3�[@����}"���M]w���$�7�����.�<���[Cq��(����͇��Z��+�&C�dAfy��|���e�*�O����pK�|�����Ls+[��s,}��"��~� �$� :y����wt�w��͓0�s��@n��. ��n!��g���X�"!�f.��cTe.��-�f�!qBt{[��Ԣ-c� /�	d�-�9���gq[�Β��amDrD�\R=8�+�B]`�����O:(YN����P.i"�7/�����pe�#��k�\n��gϩ@���h{]�;4�i�u�*�Zf��0���WB��)���TXN���>��7�نv=�H�gMm������_�A$�2d)ljL��h��1I��g �
�/�i�@���|�J�xF���>�M&��k0^D�X��b�~��+�����x��g��A���Y6T�f5��D�7=M�$H(����5yTϿ�����d=siJU%��&�1u1���{Ɣ̓��O�\<�6�WW�4��	��Ҹ��-$���ݥVy�ۊ�E@��rհ )B���K�DN��R��6�>��(��t��0!B���mFe�jB0%�d���Ts0�Wm����f���D �%��Qc�
��y!��3�(�%��'I��t����� �b���<�g]����#��W{/�����ȫA2J�҃��������i�L?�l���4/5����_Dl���$ets��GAV\�W(�%/>�B��������j��C�?���/b��8<:��������ӎ��"� ���_��7�8�f១�<`�a҇�ɤb�����Up�!����a��p�"eZi ����Xh]��WOZ6�$(5�q����$�ʕ}�~G�kt��:�������}�i�KO��U�W�'������D�͙�bܖ���0�;����RZ=�c���_D��T�r�>՛$�����
, ��܇��V�LbO.�����Z�㈮5/v�->�7+�|����v�|�11+��od�|=��'��	��������k��,�9�����_���E�6K࠶���/O��t��~5wg�S��Z����Z�<K~�Go�[B�z�~����?4���tPn�tH�c5xL=��)_�W7��c�c�ȣ�w 7�E�#	n�=�Q<�+y�U�����Nͥٙ�x����1����|u,��Q�5ʑLe�R��2�.<i��`��;�R�Gjq�p�LmwJ6AUښ��&��,�t)XNҖ�|C���.���:�A����2e�,���L�{&�(��bEC���i�*�Ȟ��N��=��y��� 	���5m�ǭU�"�5�2�O�g?d�;ѱ��jZ��)$�*F��!I+9������i����R��h�����3���/F!d2g���0e��pc�qN�̇h��w% �S5�q�{���:�a�y0�bS-*������T��z�}�Lu�����l�UG�cu�?�tz�E'L���Pk��#�4 �6�p��w�ԧ^����L������$��A1�ėI����FA�(,��@n�Pn]���%��z�g�$rSwS�ؖf$V�"&3���H�<�qH�ʊ���Y<-�s?&b�l�Z����(]��%�K$�7���������p��ڒv�L0�ɦ���[ɭ;���Z՟G�U�?^�d���"@%-�G����L���	į�L34��-�`�WN�g3�s�����7/������6��)0A��2JZ6R8VQmL�=(5����̐��ꀱwz����>+L�L�7DMa	�-�m�ʨ(q{��"���M�Ԫ�=.}���5�&�s�A�.#�Sl�t�����C�w�{�:a�lBx���J��9�Oὶ��{�]�h|.;�Z���]�wmv�� ��0טRc� ��b���{@8ѹ7��[[ȡ�r4��3 �3r����T�q��A<ө�E �����U͏�(M��n�t��c=�X�ކTO��Hnf�B�9U����
�7��ƄGY�� y7u˸���8��a��V�Z�����L��d�8Qi�(�߶%EA�b�.&12�Ǜ�|�%�@����5oG,7���q`��9�͢m3%�x���'�P
�ڬ� �yݙ���o7$�=ψ�Cy�Ճ�q�7��q
f�	P��F�
Q��\vn�Ck���%Bo��F�<�x��l]�%�  �?�;���1{$w����,[i�}c C̓y,V��z���Z�H9x��RNE� �����n+n�/4Q5�uD�m�γ�-��܊iq�	� o�,@�w��#��9�+���AZ 
[��&�e`a�
���+���b?���{��~P�d=W�M������|.��z���_�#���L�%�z1�mde�]�lf�mp�YP� ���g��ےn�����N��w�ʵ�����y$��_X�ZZ��K�(�''N=��ދ�Q��0����8���nBl���?�� Px+d?-5�T!�0[a���!�qj��}����y�������b(���=w�s�L�s�5�I���\� C�`��T'd�ީ�"���QL:
�l��*y/��{|^3a��.���O�{.1㢗Vtu-x�)3��3�L%B���1}��b�1bO���zc:^2d��6����z���?��A'�2��ȃr�qV2?��^�&�]�����И�̙Ag�H���n����P4n["� Xy���:[f��^��5;�0܇]�L�;��D�㎮W�o���]6��хN4XV��ǧ�3�Ug8��Q3�͵cԆ�h*(���勃���n�ͤ �I:3�����>�/�d��#����=��9�ٺ����x�[N��6x��Y��A.P}d2���䷽fо���ki�_ꎁG���\��ৌ�35Cfe��!��E\G*\�n�Qn5��-��O~$���"N�T�4���eԨR�yL��`$m�%����d�^gd�?�dݨ�6�/�%?��<|�0&8������-�$�^[/�nƒ[��b6s�r/]@����)�����yn0�*ʾ�{�c�6����j��[��&��`��v�C��+hH�=����+\��|d1Dk��)�Ty�e�[7���8f���i�n�x���}Kg���y����N9�h..As�%�3�-��
�c	9Z;X�uv6#�	~�S�����o�|����W�����i�5������C[�?&gFk+��*�@�ʘ:٢�9�{ K��^����F�8(ט��:/�S�B3�֭G����Ɖ������%�W�]��༶�LDcհm�~$X%ؑ��|�_�Q����!����.j��f��MA�xR��?!�b	�R�|�
�c����_�A~n�f�gǎ�l�����G����(���{��/0��;�B�u}�*B�R`eh����"&s�1K��R�D(��/7tq�X�N&W�փψ��6�XlxVHYEB    4f62     b50������z)��>�� ����r����Jnp��4:/���s޽ڂQa\�[AZ!��ʛ,t%'�R�jx�.v�l����8�f=ω<����smepub��p��v-�eH��PUs}=h<�j�h��:�qDtr��+��+��(�.6g�b��~f �7A�0
�R�xBp�x9Q5ush�*�������quʤ��WFl�����q��}۝�	��\���-\�A5��!r�X�"���n"��+�(�9��b|��Z�2�M�����N
XO�l�V��H3W�6a�$w�%����{n����X8� ��=*t<x<���ԧ���w������Zd�0�J��JN�q,�|+/ 4����O������C��������ʘ�{����su����.r�QԒ��a|b咅Raa�U�j�k���9eK�����~ǔ���#�Q��|�S�T��'�sQBڞ�sꀪ��n�#��u>�M?� �p�cAϹ�#!��y=�g��{��2���Rϧ"h֢Y�8a�P1Vxjץ�* {��m�D��S%ʸ:㎋�!׆���&�9r���s���������07&�	�!�+�q�0���P�=�}��	+J�n���UةB��GJ��T*zkt��@�!�E?�Jl�6����x��e�w����O�*�4
^�'+�٣��a�+g@(�I7�������ZQgK�͡'z�����!7�i�����ۅ���Q�/Ձ�w_�� �p��}���ܶ�X�z~y�+,�f�֔j�]C�|�=i����wS����6+nP�n�xo���"Ew��v��б7��wVo1Ljc��+�p���Y��������n�@p���oy�XL��?r �.��4��Q����L���?z��/�5����6j��L����1�Q�ܔ1퐾�.>-`�%2hu1Nu���@�l��pR��xw��c�?�������#B �rU�U���k	^y���\np�ޔ�b�>=@N�Ċ:�K�����)�I�VgC��EK�'�V5ɇ���g�vvÄ-��mQ�U���P'([�9�|�i�v��)��[ ��k[����g�o���]ؤ�6=��KF���|`�����&����0�'�+լ3��WKY�}�U5�J%��t*�x���Z������F ��3FG7
(�3��Z���:3*�s�����w�:U�$���L�[m��m뽍�wՃ�2��>]iŸ�*�RB�>��p���Ԕ�"P����CS��/���D���Uy�<��h�Z�4Ōb�^NV�(������d�;Q�R�U��a>��0u�㵢�]��^i!:��?P�N*8��t�G�
��#yg��saQ�+�e����%��%)xZ[�|�eL��U���ΠS.�cp ��rJ�(v�]���[�wE�;�֍�YT1��-���׮��!�{,4�O/�����]�"�n�_pL�W}�%��������2�I�Z�Q�@�l�@)��K}��+�������۠O&i��c�1��Z|lgRِY,_������b Θ���p�aI�e���[a�t��Z��w���G�n�b�[�ҍ�������ʜ�t��X9f�����m={h����{���y^'d�<7����ڵ���+�G�Z����?��@����gn�����<&���5���S͒��b��V�Kd�ۧ�ub����V�7J���QR�
���f�w����!����Ja<W��D'���ۭ���|���* ���t--�Ή̵�O<2=2�3m�p�>�*������3�F�������"�u��kA���Ѿ#gȆj�rS�[�G���_<����V{zIBi3�B���l����x	D��'�T,�Kֺ�V���("����=�%z�Qv�u��	��@����m�D2�^���򙅴2�����혗$wA#s1��Y��A��"��ؠM%�8�2Ϻ��ۚ ZV��A�j� �h��ڼ�
>{k��c�z��e�����^t��Ns�X�ڎͤd�V���i
j�Z"!�JZ:a?�\�%���S�5�m��o�Vl9s�Ԟ��p^6�z\�h�p/�}��줊uq4p��Wx�qM0���� |����v�a��y��V����SV�%��rN�� ����MLy�,u�J��ww��W�dx)�R��|����
}�_�4��l��D$2�|�C�5��GYRbQ'��_2�eۢ�ע46p�LiN²I��hCy�� ���xv�����Б<X��	�p�
!�V^t��yr0d��ֲH��bs�������W�
P#
�82>A��:i0��@�A_⥓R������p�2�_�!���D0����%�����N)�9�3h#Fy�$xd�X�x:F�l���h����B�lק6b:��^�Ή
>H��4=�tc χ�7�G��H�@�,�M`B�k��[q#P����"����9����5�h� o�����<�l�?��]O*;��+���xb"u���Q�O'<&�D?w���J<�U�/=3j�Aq#��`+2��������B�wN���#�-;����#L ^h+�MQ�l��?Mo?7J�u.J�N��gV�+܎�ݬr�Zw���S7`
��r˼J��d�Kg+��㥊+�";m�Cu�b��}O�G��A1����������l��%�g0X)��p��)ᾧ�]�~TH���NX�.�b��v�x����X保�
L�Ml��J���y��;����v�5����$�Tc]��RP�&�W��V4o<GR� j�< q�1JK��}������qd��P�3dS���I<������4��i,�hդ�[�}/�o6Nv