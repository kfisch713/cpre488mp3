XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��U4v�,1�ѷ�7^W��>�V�dU����*W=�=�R��$�\f�hv��S��IF�}>f<pKl����T�t�u�q1�#z�`�O�?C�����aɥNa�pb:%��Yi�76r♾�4�P��B�<i^�"q��.D���B��1LfOfB�~p�������?��\���ݼ��j��&����T�]�ʣ�q�;$�i���� JEYp3�K���N�$�J�:����g�蘄�7�l���	N�td k�ɨ�o�zu�j�%�(3���.@.��>}�K�MCx���r�k�D
�t49_.a�y-r�;r7*85���1y�5�������)ڳ�>� ���%{���;q�sir�U=(�?z�� 
�O}S��?�-�e����"Z�Тɚ��_���~o=���Q;ً��A�-9��|��t��a��6KR}Li���8�Ϫ�+�R1�MY�6)���hB��=��Í�s��G[�p���O���z�)��D�mb$C1A4o�`��g�M��_�X#�Jl�k��E�cV�����K�z	q�|��&�Fu�B�:�$^Pi��8D��F��(�Gs���D�+REwr��r�z���=��g��H�����GU�$� ���/6��!k�G��^�^��2Bs��F�H�8L��W3��+�Sȧ���Jl��5�q�� RH�C�M�|��ңELְT���\�U�o���r���4嘄�lW3�%�r�������]Y��K��K�T[�c��xݗ%��3�XlxVHYEB    5d29    1390��a'H�$HS�p��ȶr&�m�g�L����4���u��S� ��s�pL)��S��GGYٻڭ
d���n��@i�����xw�O���!Ұ�;`^��7@�(�SF�=��C�X�I��'�fK �����G���͡�0�fG�_Ǐ�W���o�ie0u^��yG�gK�kT���-�9t��q8���y���1�ꍯ���W<�;k8#�oA�z��c���D~�{�p�ۖ�롏���un�!!>J�/�����[��A�pRJ�οB����&̱���H�KC��W�z�|U}�HY�}�c�&SЬ�����&��A�X�NKfЌ��<D�6^�(�Mqؒ4����Yw����ٔ�(����lɱ=z�5�� �0�M���_y\Z��[jgU������)a*M�$�?���\~�}I�8�!���fޔ�%��v-�qM�]=~w�oJ�p��Ӽj98*��^���6�[��2*�(�^+������$;��<�$~W��H�.!~�!����2��j9����1��$�S�Y��;�:�L��@$�����n�o��ŕ�g�u��>5m,�_���zLq���r&DH����O�|f�j��t�|�Z�;��=�A*�-y������ф�oG6���Xb5t���_�eN����|_f�ҦbQ�x� ?2���?�NN.�}9�O�˹̲��/�������S$���v���.0�����.�h���4��n�#�SK�y��#��<�ˏ>�M]�ߩ���S��^y�2���39��8�#1�D�
Wu��2>�k���ltm1�/<��ܔT��z�b �.�"���Y���0���X+���7�����B�J9�Ez9d������5��i+�a%�t���4+r���HGl�њ~<�E�����VPk®����<2W����n��2:<�wknB�B�8�.�}"rc�d��@��P�O��7'�'Z$�N�x�T���������C�ؙs�E��l����#.l�<}��H���V	0�D��CV���4ӠbK�S/5���V xhi�Q�ޕ��:�dk�v뢒fVb�Q�c�x� �Q�v�.פ���O}���C��<Ӹ�f��P��"���?M$��TF�XZ ×��В[�>���X��SPפi�A�л��"��C����l��g���լf��V�f��l���? T���Qv�H�;=G���EϏ�� ?�Sc^j��Z�8��rm�g�K�����:9��\��]��_�� �1j�-h�3v��W�v�,k��k߁�8����u�������pAz@��z������4��ӹ��x[�<�%�P����9��$�ఖ���D��(�\�,���
����`�>h�Q��Ώ��z�8�Oօ��O|"ܒ?h�<}*x��ɻ��:r��t�K���$�w/�о�{7*~+�$��w�a�`�6Q7�"1
^��?:ڸ\en��Q�e{�<��[5�Y�xX4quQ��v>]QN��:s�`����tu��\��42+�Xv)p��R%,{����ө�O3�S����L��;��ڠo��Y�RXz�hq����Я3�r��a��ƶ��KԱ�a�X���~?~ l��1��r_DӀf�OHp�P�D86��5Us&�i��'��	��&����K�k��X�^�6G���<!��U��Y=��,�"*�ڵ7K�6^#dHNξ4�Pl�Y���&q7�m�5L�}��CND,��wǮu�m���u��Q���.:���L4y[����Yq���GZ�@�Z��@�SZ,�$'��G;���cxIl�����n2LrU!��A�I�Iٽ9����Ǐc���;�{U�
��`	?;ETBHQV�ڛ�d��Ӡ �q����e9tS���p^�'lrȥ�� [z�?.XR�xQh1e>ћ~��?�����/(�&~C�L��E�:�.J�l�]�%���jو��?���5���! �a�456 ���@o��b�iB��5�MJbxj0"�E�����u+5nB�����ܨj;M�9C��d?% ��q	6�0�\��������|l�J6��}Z-.X�$�!�1D�K�޼\�#��φisё���A1��Dn������g$����>�Ǡ���L���,�	;o��Ǖ<Ͻ�!�Z#$���]�x��F�?~w��Y��Z5zrR���~��IW��m	��*x�'澈|]��<�����tY��h�����H�E�Ɣا+����8�l��}�/J@��>��/��P�(�cI �����;$Y���S=�}0��Q�y0�����h�7��{�g�e�i}��ؚ�k�|��w�e�W���	J� ;��	(�$n�P
�O�?�ȼ�)ZJ�E��{�ҋ��rN�"򿤕:X�g�?����&.dƕ�D��)ēj��Iv�4 ��Ǣ}�l��ͱ;�=��#�N��{v�"	%��H?�[�0j����Q[2ZYJT��"��I\rT��PEƼ�Ǽ�\�i�J�`�]5X�	������B-"P`�eZ(���T�w
b��v���Qq)�`��'ߜ[#%`�Q��ȋ/�H��37dm%�+13��X��hk���0I���
Y��%��>0+]�Q����b�0��6I;�׀7kWŞ��� 9pPc�Y�]ch$�l��R�GI�
���[҅���ù{1��<�H�춖�4Ꮾ8I�G/�� 
{i��t/���%e�Y��-B/=�BP��d�o��x����,�[�B�&�G���AW��E�E���(��]�҃��
�������V���o�zYk.)1�G�}���_�5	��nV�`h�kn�䭋��/w$$G�����>-d����#��	��"�p�$�X�FX��-��\']<��~*�����P��H���kJ��	(��qJ$�t��G�*�������lm���\g�,q�(�X
S�%lx=�� Ʋ�c
���Ki�Ր_o7,q�n�dq���%�L��>'�S�%��M��
ٍY�Ο
!�|j�O���L���ֹ!uh��$��(��)�̋rHZQu�aA�}��J��w�b��#B"s�i��f�Ȇ�:ۀK�C��F�V���r3���B!
��r==U��
V�B1��k@�E͐4���û��)̢��B����b`	,�6t��>=r��:�~��J-~�@�`�R���:��w�`w�E��h|��[�6�Ҹ�G2fo�Rk�?����]+|g��otV�M.��}�ҥ{oYZ�'&zhPP��?T߼��?I1�θZ}�����T�ɑ̇����}2�_��o�uw�$m�����Pq��p�6�'?�!�&���]\ ��~�	�	�y1��<!���>��f������}/Ix(�Ȋ��������5���c�`�E�»z�d_��28��R�kFO�����\�s��I��<�-��s�q��Uu��)%^�	��1$|g�O��o�,�y�/��R^��_��✄�]��!.bvNj���hqZ��F�mP�l�}瞌���{a�"P���'rؔ?���K	�Dk��\i���Jߐ�gF�T2�Z�.9��o!�p�v=�
��܆�x����q���]�E)p�_ˁ�&����A�>_O��m�jB�"�9���\ǂ�%j���k̗TU�_�'}����}��%ַ2Ո]�X��*�L�k=�nw[
������h@=�,�ӧ��@L�(� C�7��_��c��[-C47��C+���H���]��C�3x�^�,��<DN�V��o�arT�� ߛ	���.-2:��?�e�"���۱�Х����ߡ�U6`ڃj*��'4B�(���$�S_��9`���l�O�'���8�-h3l&��G��F��L��-qB!]�ҏ�zn�1���_-�dc�YQ��y ��?!�8OџPn��_�k���0؃��u�^�t�\�J�����4��zj��݉Fܤ��p�J#U�4���F�&��Hb� �C>�c�P ص���h�p�3�|V�������1q>GA|��P��8�	�%>72�[�މ"IW�q?����6`*U<���~Y�/�]��3H��܃>����db{%�i�9�('�%4��1����2m��v�g@�s"f� {Q&���5�X�`U�F$7���E�f0�5�s��t2�lg/��bB�?z+os�;i�kq".�E����H2 ��`ڥ�oe�N4�@h0�A�'�ꥥ�ފ��C����!�T��YYe��ƛY��������ö�z�� ��@�ܭ�Q�i�Lpt��ǹ�tt�,zEMS����wi}LT/��UR����D��ӽ���}�p��V�L��{ˎ��|��e
\��[�Up�ga)4nL�@e�H�;e
�s�Y�^Z!	���B����5�:�pZ���(�dc���֨ę�)N���Q��=ކ�����\ �Y���b:x���x
cMnR���u����Ջ��>����k%��۲����n�=�DHL���ӊ�f��h|�\`&0$���\��]�kxw���0�d<�����:1f]���t��C����ڟ���I��QƁ�f7�$W�W���ó�:�aZC���c�v��sE��<�l�+���!ӹa�O���L	�����E:9��;
������'U��1j�A+�8Dѡ$�i�]G�i�X.@0���s����3𨆂Āgnh*
�p9�]r]h>]p����� v+幍~���oծ�%o�zD�a����`�n���BH]��Za�*�
7O��V�	�$�-SH�{���Hz%�W���=��g��R�>�����$�>�� 遌bb�Z�IG���������×��!�A~�$9�i�M mΓ��