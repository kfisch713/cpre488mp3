XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��ep49AY}�ik����a�����H�, ����տ�놣:ʛ�kZ�&�jk�b��v������<�0�d-�K,�q��4�?��g'���9����������gM�b��o�N錰��\�j8�aA�tM�K���=�����=(w?�:򴟣�%$��T�w�,\���$��2��|B�u��W��b�%�V��ɔT#���-?�oT�[�)�W��=��b�F���l�{���u���h�+�2o�mލZWG��|�$�6^?$V�BѪ����4�KCn>k�?8K�-��}�L�-ܦ�"@��-�6�M�$��|�z�ӡ-���Yy�Ӣ#
3�?Y�AA����o5�7J�Ad������u;�V�B��Җn^�r':�R>�k��SD��lz@DIr��߫�!|-=�ӝ6�p�=�P�4���bfרQ g�^�	1��i:�S�a*���>���:��G��Y�ύh�71��V��L����S��l�I0=:E���=�!�>�?�F㰜|a��e�z��5�q8*�����K�� La,%v|�ds���]�)8����~oZA#��_�G۸�e4��9JL���?�{�ҳ���K 6�zf �f��e���*��Q�q:�s"�9Uh77&�U��n�1�1a����
���k	���-�# Y$v�s"�+ʹ����Hl�2��M����{�j��!�	���'��N�U�3L DK�<������h!g�ٶ�$�	i�qԃBJx8XlxVHYEB    2b75     cd0�J�M������P�����m{����O�c�GMH_`�L�>S�LY������d �s�|�M,S�L���3��3P=
�ht@�	�(�F	�f ��@Ȫ��&�Q�qߍr�1��2���~��yT�W�@P��	�2�~��W
�������r�9 v��I~��dii~��a\���"ݦ���"�rr�dմ��F��s�![��-
�ʚ���.S$)u<��Oܡ�5�-����?#e���r��q���� p��U��zk䲅��d�{��&�t��b�Kɐh�F{7�c��a�r��=�v����Uiߚ�V	�,���Ó�g�_��a��q������̳%kF��c�r�Zbg�^��L��W��c�4�3Z�{��Me�3Z�|�4�ȾZGs�[��D�)M˞&�#|[3���uq?���Ctb�F��Z�82|�`2�:�*��/�"����E��/�v�U��YBJ������a�B��.X�$H2P�}q׌�W�4��)]����=�Vc9��ҴxwS�({�*7����*ũI��\�>9(��㭙��,�X�&� ��&JPM��4��*�!j��9o�
wf4+C���yl��u8X ��Zrw%��3��GK�������0Gt�\L|~���������%*�6���qvx�V�k�� }_�q��m�Q��y��b�H:ASڒņ��!�@,Z H��p(���T���8�눏MqG0**$�>� �R��81�
ԟ�EC��w79V�V���ʁ38$U������ʑ�)�܀�����r�oK읮�Z�{�A]�3�Șf[K����p-zb����E�W(��L
�@�.B�T6�2I1E� L�>Q��!�C��c���ɬ��Ct�	���H%��B�J$F��
ܝ�t9���-����X��� W���&�d�����ɚ]%��JB?a�����L^�.~yg_�4ߎ��s���J��%�o����8~B,U�/�"�)�w��D&��-��di�6Xݯ���� ��_�\1Fާ�E!ceد��o��2����/���Ƞ��ae;(��j��Œ�����%�L�p�˓�H����o�����=�*2�7ܠ��4gtƠ�V2鹮��_�쌺L�HO(���3�����G�EVL杨(ZoD����5��W�}�;g~"~�Q�����d�,��4Y�=c��f�� ��{Vn�ՉY�܂�f�Pc��91 T����u^!�t�ǡ�>�Kˮ�E��Y 2R���
�۔0g"�A�&rzf��wWmN�vٌ/^ ���q�T��1��L�.(;��	w}+�tI��c��s�~<�=	�=�p�p�O�z���B�(�l��)��oq�y��v^ny&z��a�.�o��' �J}��a����m��n*l��Ř�)T��ؑ��健��������Xijqt�����g�.@�ݶ��m�{�@��B�.E3��hx#=�3��"���]`���E[f){�8&wy��B�mLu_-�6�+�i����ʈV߰�b�>1� ����EX������yf�P��bS�zr��4tb�		a�����HM��1��	��Ԡ�I�qO����|3Y>K�O;i^�����ǾE�5n5�|���O�Iߢ�Ko��m\y�_�XU��dt�4��1�^�y��6�p����x囹 q�4�����=:fi?-1F��<���a-D{��~�LTf��Z*r�B�s����~'��~l�4�F�,e�1n��Y;G(X8���5���� ���1O&�OSC��[M�Z����E��/��>�w�W���Q��<e�	�U�^���>:�ejS�|���U�e�i!�6��ƪ���/��e]5�/I}�����߉���x�Y"�3���uw����fأ��g�#��ˍ���W����o��	��.RGǭ��E��,ڈĨ�Ga.������4$S3�=�U��օ<�03T��P�2��Y�h��Nh�\VH5X�n��~���W8�9hy8�N�?p]-��\u�(��_��!Fw�+Ѯ'T��Fg��Ŵ>|�A�2�Z��'=p����	m>n��Q�@	�aw�y?��1�pfD�"��~\�n�hm�赥g�N�M��I+euI�ܨJ
/�_<��$c���G�-�~�Z>��hsD.��Q*�O4�k2���3o���s̙�&�^h{&9�J]�%tW�-5����ˍ=z�ˢ�_@&�34���ZZJn>���D���AM�{����T��a�1]���F��o��c(7hwSR"GNe����=��	����ڠ�8���!��,��1��z�>t��j�a�`dO��㝒�U�ǅM��)���+&�����!�#�E���
7�zk��Ԍ�qꤙ�vj�4�eg��Q�����)���m���^W�#�/fP��|E$�P�t�)+#�@ C/� <C~�9��d�	��B~�(���$w�����ڌ��P�~��%N%�@~��9���5��a��%�XX��"�'M���q~,K|nո���s$���e��_YF��Ǭ�\y��Y*	Hu�ʵ�ةP�G�o,���A��C�l%�p�� B������6ͤei�$�d��F�[N�} ��/��ո��榿*D�\��&b۸���hҕ+�ዤ-޵�_QN�Y�V�	*�M��ǐ���n۔��f(A7'CE��YL͹��~�S��6[�#^�S�� MΠ�=�(DG$�����64��u��1L��)���`�7<��h�P�x}QJ{��;_��n�@�M�G���F�A���ڕ��%-r����jR��`�^�,�"[��s��>s��"0�l!���Ä�,�5x Koyr�C3�~ʚo�����h����yqtU3Hmm� "]v�@E�m�WNR��a��lF������}�z��%>m��2�#,�Nx+�E�[��mi7��y��i�.���d�5L#}+X.0lU���"�hn��>~~H%�B�T�"�� �c6�ed��J~	��rV?��e�yM��jZ���k�j�`��	�CX%��Qq�HP@��Nkg���3�$��y���^�1A�ȍ�(@:�S=Q�?������@E�G5O���P�D���)��pq���FI�}W>g����G+�y�;8�I ��|�o���͙4��YP����3p@�7�5��tRv�J�w��d�0Oz��