XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���R��`�N���d�sF��V2&`�W�n��������F(� )�����
K�0��/�4+  v�9%��b�}mf��/��+5�Fk�]��z{�<�@��Fj����Z욧�!'K|3sB���=���D�BN ���t�Z���98�9�٠7J�N��x�j���R������	�Y������[�U��j�Dn��ާ�!�;���+'}��6u��<����n�&����cfA ��ڢ��.y$/��t7d�0	�?������Q�0���])��w$kw��A��1+���@��d%��#�(��xЈI�ח�z\v�wmr��y���q�+U'�P�'��x�lILb���Ifx��������H�>�����"4T&9���7�W��?@�i����k�M��h�G\Q�E�9h�Z���H7��g��;Eb̦���s*;��g�m?�X"��e��L6�
�Bư۝�.W�n0����#�4���g�=�h��lf�a�B^9�|�_�
5��-�8!�sH;�F�b�c��'���4ۗ'�*���� #zNF�����ޗ�	S0�߁dsb�!m!�;0���vЎ�\���ΰ��7��T��ku�q�� 1��4LP��7��ڏ�*���Y>Kd�'C{�Գg��}j�
VSZdL��k?N�]��	����ފe��Uߟ�>�C�lC%�2Y7�M����){dΪ�_�P!YҦ�.!���M�9����|�Ms�m]��#�yV�XlxVHYEB    3d1e     fa0T2�� �
+C��w�F�W^�ͣ���wM�mq��7`���̒hZZn1���ǐ8�o)��3�>����;���ǲ#������<��QY��$�a�)�{(!	>�}� ��C�B�w��J]���+$�B�yn4��Mjw6���:�tz�עz��о�Ɣ��-ۚ�~��Wb�S�Qˮ���c��=v�CG`��٭]��ƈ:2��+_���*2F?0���p�~����P߷�bN��#"搅0�|�bo�>i�p�ϲ���kY�F�S����Ɓ��cwF���`�]�Xe
�����7{E�� d����+��iJ���:��E:�]S��?q�M��FqD�!�KE�$���3U11��Y:�:U8��2z�*÷�����T�-�I�� Z'����{�)���Z41��ʿp��{f�
�_�Z���B ������ �3��쐍8���-��;>L�;���{Ϊ|҇]�W�ߊ�`�b�GnI��RA�
�+C��5I$�~�ShHv��0(H���|jv��<�ɿ���I��K妭����� �w��i�̣��4�Π����3��s�,�GhH��5ꭐX��� �&|
c���[�/rؓ`��qSB$�Dtײ��+�c��
�ʨ(A����՗"�a����f�ӎϙ#����@qJ�60DR�}a���=���=��'��+;qZ���6mxY�ڭ�
"��,�����w���`�y�	�:��[<�2�+}�a��©�+{��{�V�ۧ!�;S1e�� z�!�S�%h��"N|���P����M����]l;��Lf����,�7'\�h�j61����|8��wkC��K�-f�?'AbP��iڔ~QEٯy�7x���r2~&YJ
H���7Fj;����I�{�Ǹ����L���r�lű�3!,���
7K�2�y��%u�#P��I��0�$F2{n���7D[§����~vp��SYl�Z���&F6 �}3��j~��GTz��c�5����x�1D�L�-�	Ǒ�|�"n�uu�׎a�MPHi�% 	j�֣��2W
yyK����$R��u����Дi�Cr�|r��#*٢��a�1Ą �'dV24��~\%���I8͐<�J�)��	�(-߉z����I�I8M���,4IB��E(��\�L\,�2j���l��_����]��"m�
{\ܑ�4	���BV����c�.���X�]Z�pF\�b5P5�A�'o�B�DD����Rh�b����-;!tp���0v[��?�s�qc��f��3�vܕ'y�4wFpW����9
�H(]��͓<%���25�;#�P�̴R���H����Z(���K���HQa�؜�١�fi|5錼�ZK�L��x��aƟn��{���@���"��R@O���i�+:r�����P��?Lݗ��d�D���g:�D�Vc\@�8�V&���!c�qFm�{-MḙH?��A%��B�x��?q'�����c�i��\?5n�Q����7��oC�j
�������WB�9��M�Y�wt�&�w/�{��|U��!v�֛QlZ�ä^��{��a���R{ec�X���(y�'�u�/�b���0e�m&Ճ���O-�����Ͻ7:{����O~����@��>~?�����O���l�R��b���L\qi`�k�yk,�*�C���i����=Z���k;��W��Ϝ��A^��[�v�	����F@��Q��}ڢoh�w���d�EޒB���C�}	�mzҸ�-�/��(��J!�.�t�w�,:y[��$�����vf#5��P����zq�P�r�C8SFu�'ۑx�!����x�ǡG!�r��U��FIY����7�x�H�ܞ��œw}�W� ��;��)�a"�7�I���gdk��������?sҟ[=���jm��ɕ�KO���v��d��Wc�&~��B�^�Bá�Պ�b=B������c�!CG���Ÿ��>�X��eM7'-��[��#T�D�Q55�ݖ��S�U2�4Md޸�˹z? �{��!.�~���Xě��4�40�%d�N��2� +�s�i�DWǽ��h��C�W��#wb���G�H"(wӮ�sB���@#I'��:�~m`�dr�|Y����'Fs��XQ�C�_C0a� �3]�!}<��C���nTtX@x���_�~�� ��{d��
1.����+0�L��q��F�B>Fo]��xP3n]e������#f� 1<j�����*�)�%I�/e��@#0�ޫU��  bg�<A��򆍚���~!c{6jF�$zv�L�l� � ��y`/�N�	��m���I�![ jW��g&X�YxXn��ȓ�!�0��0rI�p��*��6��0�s�d��.+�f���2$<em�B���P�O6�X
 �`Yp#}�')/w��{|G���_Éi�~��lyǭM�_ܫ�o��Z��`��Uq�)23L_�=������B�R��8�K�]K����t�ӥa�Q*B,@�2����n��GQ�ah�6���F�C�Y�E�6Gx(,�!R[�7���)�ʃ��E�Kb|��?~sh��h�0�%�X�t��	K�H��M� �~�J�0�����ܸ$�f�c��&a�
�MS�Q�	GY�4K(��Y�"��uB�[)� �P/�7+[o|�N[F0bB��� T?�@w���+U�&��ׁ�����]U��r�S����5 .�9���3�(��ڬ��������P���)G�Ч�8>Iв�{]At��ɪ�om[� ����-'��U�+�rmenj.�TS���\YVF"f,?�CS�[�����ԋ���ŹAm(UVj�#u_�~�H���3s�Dx$�9��b�}P|GO�1�ظ�?�M*���@��!8.�k��ŕ�88���;-�VJWos����:d3�V��]|�#�J$_��ٔ�5��#R�J���׸�Q�/���s��~�Qޅڻ��M4B��x��5�{/������ �nqB��Cyg�#�=�u�]��i�x4r3��ԛy)��'���`@v���3��^�X�v9y�IjR�w��,���S/�u�n� �}�8�J�NY�aK��R +EsUNsH1;��F���Q��W]-��4��A�x+��F���B����q���ߔxq8��z*ϒ�\}KO�����q,�
�rD����(�R�S���!p�9%��J����~�)7������	�SBr{yu��3�6sd��. �
*4��3\���*��˧���:���k�N�e�+{S·a@��tk�C۩�/KO���?"�>t_a��  cm��Y�u���o��c 0�Dْ}kL�j�"�"^�g��D˛�G�H�K�-��N�)���"8
&s{������w�g28t�'aF]�}9V��L�t�L��d��3��|Vd�H(MiS��u���\K��gi�g�{1�����,�]��Q��������F~]v�+ �����ҵ�"��N�=G�i���¯S�"F��fR=N${�Y��҂,u�Q�=qRK�جbMٌQ���2o`
u/R���Ѕ��UXr��3!��3�QDˏWR�(��ǣ��$=����"��h}d��5{�ݞ�ʔ�Ou���,�L׊F����ؒxy�]�Q1Z!�-��3z4���5Z�VF1?�N�k^�M�(�廵� ���7x�,�����6��_+�ھ�+6�po�?z���c�D��4w'�qb�!�~�t"QV�"����j��-��#�5i-��sÚ�T�N��d��-~[h������5@.��F.��f�u��^�9�{AE�'c�dΆꐖ����U���JO�bm�9}�9�ryDBI�����N;*�t�F43�PŭC�W�[�6��lm�P�F<Q����gb ~x�a'{��