XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Bg���nm$�J�R�'?��w��d��/��f�a�	B���"�������L(��/��MY�ٟ,K2+ٜ��U����Mn�?��;���Z�M=;G�Q�"����Kq5L��g�x׊��W��/�E�f��"�����cUkcO�����/eHW�7��^�5X��]"z��Rk�|>�����$��TGy�D%�n��(�����-�2Axfκ�e9�b~v���WQ;+(nn��v�QћF9����$�Ï&5��W�$<�8�X��{7��[9�v���uƁv�Z�J/��|Fqr!&�K��m���x��K�=Tz��j-��y���5�_K����8���;|#��+3��)A�ߒ}9q�����k�o���a�U�Ѹ��5	է��_:�}H�P������,�ƻ�Cz�U-���k,���څL�j����%n"B�p-�х*^Ѱ��[�٬f+`�vL��^�%�~����"P],#϶
�R7�f�:Ɣ[��z��n���A��u-�U��4 ����ѓRF��u�?QƁM����我������ k9^n�,pE�C��*gW�DvsbY��Uqúڳ�y[�#�q�[�h�}�g�O2(�X��G��Z�J�D�)61��جS�zO���3T�cvO�$��t�����4^p	��&.R��k�&�g;YN&�Y�$7K��4�`6�!�QW7���2���_S ���/�6jg(h��t�MY4K���%nj�P��^���XlxVHYEB    6315    1790��bM
_Qmȴ%�[6=�,�r�����:,V��J�g��$[�"4�_g}�����GT�F(B�ul�ۻڼ���C-C�L��&*;$�t�D~�u���W����Y�p��v�d"��g�2�/W�4����f�\��?��]Gq�Z��۩vzVڻk�B-�u�B9"����� 3#�l�PL��1�ؽGX˛��r�iT�͓��m�t��E�%/m��7��Y���S�^\�HI���=��I,rOU���,Mz�!=A�3��6���i�pr2On����\��պ�Wxf?6"6?��d��ʍ��B�T�|y9鋞{��z�}�$���LT�Lb��#)����	E����];#�4�q���wK>�p�|��6Hf�=��U2�Zǈ�u������o��F��wh�o���^�����U(a&c�fX��J��Q(�Ԇ<Ű��ľ�'���� �\2E%'A�^9�oVK��.��?���G������]s�SҒ,:�E�3�rh�l�=�߂�Y�8�}�_�����9��1m�����|\8�Bw�ݵ���1�:S�w1f�=n{~��~ﰼ;d߯�q���`�-M��7Vׁ�_�H���Ng'���ӯZ�k��<�� ^��G�C�WC����w�':�,P�;wB�"���m��=J�|�rf�Q���q���5���qqH�S�hUDW4,elx�H��]I�2���}���+8�ȼ�>��n��d�1௒F!'N�A�M�1{� ������X�! ��V#Z�:}V����;<�2�~�`r@�_J�XwrC��6
ߺ������7�P��Bb��;�"V�﷩����*#
?rMޙ������)���.� �5��&��c��٩r��]%�ߧ�㽽�'爉�I�;�l�k���B�X�������"���D��X'��&a&{u�|!݅ ��f{KS���JR�t��H�������b�^6<��oH#�>ɿ
@�m~p-�8��v+2�ZiW�NWi���>?��(/��JI��W��V�i���~x�Ɠ7���(UA44{�͍}�J����ڞƙu����v��#gr�a=\f/�
�3�r��<ҭE�{��^w�j��̺��0�m���7̰9���޵���Q�M���f�bm�8�P��5���-A��"��219�h<}�~W�����B�=X(�h���Aj�T =�X�4���0�����F��硥(�ʆ4�����D^��է�$в&��?�@q7����-Qu��}wx�Y�m9�k��">R \+Q�2��.O^��=���^ͩiE��h���[���D�b��B��:�q�j��9:畠���CJ%��R'�8Jb��bm�q�a�{���Ч����@����(�����Ϗ�Ӆ�ڃ�p`8Γq֩��-�<�n;��:��� �	еD�pw��'zNG��Pc���{���r�����>NYr�Ц�v{h7�I<EV0X]�]&��Ӫ]�H��Lo?�3�B��_�q'f<B�gҾ��ޣ�t�VR��Vj��X�Cx�dd��g������jl���-Kw;��>�+�o� ���ψ���j6��P{ iX����֑g�>�Frv��ų
��'d��I�t�-9H^���ei����o�#���H�]��%�\�nh�P�M�N	`HK�H��U�BS��S1h��Jor�j���JB�: �co�z 0HZ�|�5�w��ϕ`���uT���b�W�Q�V��5��-.����\(����@���_�����@6�,�x��o�����6�p/n�[0��I�l\=��B�q=��L�k��'IS�~��o�_�dBP����>�y�]Dc�.���_~���E4,���j��]�Τ�,�ysoё��h�jCdY��f6�����Ϡ��"@��>,�^"Mh,AQ���RX����c�h��1����I��xK�Ur�l�Ј����
��I��jz���Ù\�� �I7��6~��(��PQlNvOs�o�6e�Ӳ<Đs(�E���[N!nĎ�J'�Y�n�q�ӧ��[�Xi]��Γ��<�Ǘ�J	�f5�\^,������q�#�A�~������it`�+p ���cƗ�2e�dߓ ;� �g8�S"%W.L�`��t�bx����^h��V����D���z&�T��3�'���}���A(��sV��R#6��0����|����|7@���-�y���Ԝ�5�z��49L3L__qsJ�P�B�j���
��7
B#���A����OE�YC��"���ͮ(D����7P�q齃6���k����@�K��e���j�^Oz���	϶�K����-�����2�lS�}�F�<{������ ЉR�/�X�rc_u�ڇ󛩖�(uSA^iZ;Gs�Io�B��Y����#Cݹ��f�?��J�'�-a��`'{�Q��Ʋʒ�����q(�ʳ�˾q�Uڢ�����jE"'��=��ꈢwA��"�%`)�?4�zVU1BX_{E5Wx�\(e^�'��~�%M���B��?7��g���+�+A����V����H�8*A��O��v��Xk �,�/��d"�?Y�C}2��#JT�d_p�l����d�m =�tu/��MQ)�]n�3��%W� �!��oG�n#;���L���q�enNpF��	�а0v����^5\\<��"��4ub!�!e\����c��_�1�od�2$7i�b]T��R��,��&䜓�jD��&�u���vV��5�NhL#�V8�igF!Ԏ�ȧv�p�Rr�Y��Ue�ח��+��?�]���0Z7Յ��yrf��Ov���X~=[�'���v1���x�ڷi�A�	M$@&�:����/7���m�L�C�2+�Ij ��I�Z��I��6%��s]3%(N:�*m�k�7g��IqT��F�ir�&�{Pї�i,����8�����ۆd�N2�9��ݔ6}�
`>�����>�)�&��C����=�ҾC�H{�����;p|@�\Zk�?(����ԇCŊ��h_I{ӆ���$�ދ}v�����1���4��p��$�)�x3n��<����sH��������z}&������]�����W�MgN�t	b^�t�ha�� �Ev��\ޙ�>@˕��2��H*;��0�:@H��E�]k�xQۻGi��t�K�5L��� �~�<;������RPw��H��R���	XM�]}�A�5Sj�K\�T�EBw��׳3��0wK�.�+����oz��ůD��l����&�B �7`��W�g;*�~�'j��X�h�W4+�.Pd�0w��f�����s���CM����Q�FQP���e���M�d`W[h��/%T�;cװeܹ�y�A�<b��w)8OɇU �F�a�t�E��֟�YZ�ۆL��~Y^����ЕX��X
�6s�|�`�w��3q�[��V� �t��l������lJF۫�ky�A/�2;��=���e0\�x��<	/�:�S@��:蒦���0*st�s^6zr셒��V�M��U����Y���oÉ�z�6�E/
��N���9�����j	q�#����g0k�G��������eQP�vT����4�ʟ�a���H?�$���}���]�y��86o'59��o�<FXF���*1��r�?�`�Pi�{b������܆���aaF�K�3��T�Mi�o�3f��A�V�`�>�?��w�`��R)5� 1s%O��ۋ˛��%M����E��j�ޥ���L�(�_��]� �#��|pD�4q^���/��ZR����6JBP� �Y�>�`2�ӕc�9�yk����s�Wĕ�� �/ў]��;�ۘ5�	aU�A�Q3�O���Hw{�������<%�!�����2���v��62=bV�V�M"�W�g"�Ή@:��2F?(���b�_�y�p��ty�E�*>e��<��d$ -C�;��oĥ�߂=v�$�9�ǵ�#ϋ�����n^3�"$�gM��[�IA�����J��W�?�H���H\7�B�_���ⲋj����5����J0cZXv'-�"{Ȳ����č���5u:�p "	st��� �T��]Y����g�#��;Ӫ��CH1��-Xi��w�i:�|�Ѕ���"� �Z>"6l����Ǩ�M#y��ٓ�z��ژB\�_������"�^��b��+%B����)A#Ol���|W�V�_3���˧�?��:�����| ���טT�Ъe��$4Zl m6O�����.Y��/�JW�c�� �+�6��z0�%��4�~H[ ~O�醇��d�YUT� SR�1�zB���*T���My���2������H���W`�53���xyNh��Hp���0�|:7;���0�dys鵬��$E�V���]3�H��0�}��:��zƺF������XG�6���Zr�*�Q+3�]��go�`�T�k>��Ӟ+�KJޢ���^���'����4�FO5CJޡ�d�{�}5�#y��bj��Z��O}*��bl�YȃU�����h1�%n�H�^�;�D[��Z����D�B���$�Wl7�q��Ʋ0b�`du��ޙ��ֿ"����g9��M 6L�(����kЪd0s��\��}/�6��JS7�^$��Ԓ�R\>�9��Vo�A��Wv�㽑B?Y)�WZ��G��}��W5��E�aTX�Ė�ٓ���:G��gZp�y.�q���<���{x���q|�1N��^E}�+o���>��T���[5����wp�լ�巀��H_��*����b녫�r��(�y��i����h�	���/��Z�y�#����� �N^Z4i�/�7l���G]��ъ�-�~/�c��}p&��KS��ͯ^/iJ�����'�]Ɵ+�*�EN�q�:�UFI�];N���60{[����.�����@��Ɠ�Ƽ�mw }R���R*�ѩ	�)7x!^�H}�{�Ȑ�u��.IM���.y���69|8�AHȩ��G�@�P:f������Ԟοt��4���R1��a�IY$�m���*T��m�/S�'C���%���+��1�=��&���WJ��&��=O�yÂ��" �&>k�i��.���ΥJ�f�Y�]g�21����2.ہ���=�}U=RѬ�z��!h<7������C���r!��C�%ZI��$�2T�hi�!�� 1}D�/=��Z��6?�H��^�k/K �EF���!A#�5��n/�(��I)c ���ԧ��@F{ xz}����I���$����X~L��I��sɃs�r�Ի�P�<J��~`�l��m\��aʀF9��L��O�ֳ3��h�TE�� =���B�QZ�ʜ�푂�K�b����J����K��.OJINCȱQKC-�/����E_��8���٬"ut����YC�!P�hE��.IA�K/p����F��6��G�Q�:%�Y��/�6�HG�_}6��i���$lEYx�	��A��E+i�Q	|��W��	<o~���
��O|�9~�)��X&�Z�E�D>�O��)����"杕��۽�DϮ1��0�A[F|�
P�?�ے��.��V{^�x�HTa�'�����`�>�����*�̕�0���N-�.��`ޚڜ8�	���j��e��C*�Ú=����N�7�+\�%;U���'q�J��{3aQ����<���s����mqp��+{5?��%R�}��Y���d�Q<̓��p��.����ߨ��L%L��c�wL�v��)��o%Ԩ\4�����zf�׾�����d�e�'P�;�<��s�$���D�I���Tֺ�c�Zq)�FR2�q?(���e�{� �`��l�$�"]�]i@ܥ[5v�SdUқ�3��X�P��NO"�L`��/nC�P�J�`"yw[Q]����+P�"X�E$�N���4�q.?`�ԉ����n~p=dpi�#�Xy�7��