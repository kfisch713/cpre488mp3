XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Kr��X�$ꭷ��Nr9n%H�Q[�쫝 ۼ�jdZ+��	ZH��?�t}_�|o��'���˗|�2�<������Y4#�X��Pr��(Ų�>󅏢��ߞ~���ղ���j�v��s�䗈�gI����s��e38���2���m���i�s�8@#x�X|��}�����������y!�n�~C�F�󚁶�6K��I��P EĢ��f��Id�P0��φ����x��v��:.-��ە��}X��>���P�v�Z�sַq���p%��fA�$ߠ{�:�=x#����~�TM�`�lU���l$�2�Ut�M����ֳ�j�:�k�U��7��L�`��.��,��0
M��ۍ�I��X�j�3!; rҟ��y��q�2�P��#s�Ia���/�5�VE�S��/��Ś2$3������\��XE��z����F]|�7:ׁ�g��G�����-��E��vT܂<�|��`')�QQ׈}t�Px/:fR��!����Cdi�ڱ>���2Y��e%�O�V@?��ݺ]�\�*���nV�د<���^�r+P��F����1�g��=��H�l�*�;D��e3ރ"�mZ���<@"��q�`y"r�W�j�҂��ݘa���S)��� ��tPkº��>�rҍi�t�"j��Z?3m��Ŝh~w�[��Gy�����(�a!X^ �85>��gWcW�3Z��&�35�(�'x��EK�ί�,�r�9�p����f�{[XlxVHYEB    1a2e     8b0��Z�bV��~��<�HIXP0��Ȫ��?b�߂�ɑ�W�O�,N�ԝ�N/ͼ5��������Q�z��m�"G�/��a����������~���|^*�g�3���E�w��w'�x܍���֤�+�N� �����<b�E]{ݑ��j���T�������s=#3�g�l ���	}d���uT���>���@�}���	i`�߾�)"�jr�V�z�aNlL�+o�B�Yo&2T&�2�o?Y��Ի~~�"O����X'`�7���_,�}�Y}K���;}��;���ܚ�ƾت"��]��G7�п�m*�ٱ!G�t�:|��ق��wJ�V0��V?R���k� ��K�U���)�E��eCp�z"h�"q.� +�	�L5����`B`��gW���ǐ����xU /r���}>�r� �N�����M��8�?����W��wl�WBx����R:ڨDϛju��jq.A�֥e�S��I,�f^����W*�$g�h�ּ6؇'�E/:0P�e5�,0)_B۞�4 �BK�og�\3�ETZe�[���Űc�R�k#�����ׂ�xV���E�s�.�'Dr\޼zOj9�Y�q2�.��Y����ȣ��Ҫ������},�dZ�O�W9u��A�5.���c��S}3���"�K�ʅn1�~��q�)��cd�9����g����|�h�]x�D�O�*�P�f4&~g��0�n�
۲	�]�W��_	��d��+٣�	K2����"htD.�21N�˸���!� 8�� l���w;�����\'���]5������m$�r�ܙ�H8MV~��j�؜�LEm}�PsO!48w�fbD��P>��N�--/�����]<^R��t�7'�?�9\$�-}!�%���Y��h貼�����L��(H1���ߕ#��.��o���M6��GkP6I Ĉ�)����������W�<�korSb�`f�U��=fL��L��CwJ��ύ8��W� �G<q����p�j�f�f܈t�H���o���FtW2e,����M#ݰ�{`'�37��N6��Dgް��N����.��@�;�r�V���b��e��h��`��ژ)#Ko����]�$-_?�����SIM�h���a���ɱ��1�≣b][v/%�۩a�W�{_�Q�M۲4qSM�"]I�W!����$d���PP>>�������B��cKǔ����<� ��,�=��
�*�gb�:�41Ya�l��O�E�����]�]�>����G�^$N.��'MĶG_�p�m��u���蠥��p�&�V��?G�	=�G"v?� `E�t_-��+8�KA5�`|�ȵ@߀��"f��l��0g�8[����Γ��?����˴���@�3�;�~�jf,�)��֤��u��I���]�A�88���]Q�4��n*���B���`�m�P]�F!���í���ʍĄ ��)Fg`�AG(�x��S1�l��0?k���̇������<���n<�*�@Hv��<�i���0=?|�X�H��08�%�>� �/g)mX��9a{�l��NB�����'4�]/�ت�c�bY~}v��1@�(�]igrr��i(f��sW���<@�!�Y�ރ2ӞcӇuF0IX��w��L^�Wa����\���<
m3�Ԟ��>�:��9tp%yd���U{V��,�!��ǊI���a@�C�ƭ�l��h�Bp#U$�v�noH
/j�_�ogz�R"�yK-ّ��aL8�$�]b�o@��sR��PXY�hilpf��.��0z�V���>2O���G��c�	��%h�.1��~��D[s-sU8NM0�!N�/�����S���y�O�;3՚Z�Ϛn���_�n��=�D�H0���˸��cb�)t�M+L��?8��z�􇀰������kg��K_jc�}E%�����傝�<paß7���Ei�3:���"p� �2���l����$�K@#��`��vӈ�p�ÿzSF� �������[�M����8Z߱��c�'�ۋs�z
�W�J�s��gA�8���|1�_�I��]�9= ;�o<�q�D�fJ��z���8�:!���ۥ�g�U�u��3�l(�,w�B�����h��)�<�/��n�*Mպd\[�!8�* �@��Uu TK�
���r#�
�TЦ��