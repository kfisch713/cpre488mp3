XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������mn�n:�N�M�"Gۢd�o�zU�;_����6��p���Rn��L�]��U(���/ԣ�2�o�����9�BI,����ͻc�B��ձ�3�1�WPe�X^�80t%~��Qw9��W�����Ԯ��]�	"붐qW�?�N1MO� ����x��Df0��O�+�x�ȾG��c6�e��e�>�/~�+_��/XJ'��.Cf�]�4�w2� 4Z��Wz����w� CZ*����a�����R�o4���X��7�Ц�F:��s���2ECd�}YJ�h%��Q�D1&*��3tMl�`2�S������|#�=H��� Gf�2��[���B�;A���	�J��|�#���W��)��TҸ,�'H�?
o&�����ƻ��s�>�5�uEP�1N��I��fl�:���?�*���S�����Z�m��2�����-X�/N���U|i`���QȒ���^�x�Gc%ǒ�|wr���E֛PA�F��;	<�&]�:x�����
�V+���$�/�<�͛�Η����ͤ�p���!����A�����趚��:bV�/�2�8	5/�����!�"�����K��Zv���|��S��q���2�2�`O���"k;�����v�8̊��>!����$X��JK�ac�C�߀��^�bΔWH8yCؠIܕ���#�)�{r�%.gFDg&���,a+WB���G�3��R2�}�ax�����f���enAD�t����/�'}7$�:0��zXlxVHYEB    17d8     890�����`���q�e�A����6B$��[p%9�7��̏JY(벫�Vg-k���uF_�1;���^�cM-G̏i7!����8�B\r���A�?�	s��gauU�K��8��Ik�U���0K�������Q�>�*24v����o�5ڤ�`;��:� �����Y ��(�N�^C�K3��˿�O��P�J�U�)����c�Z���-����y�
4/R	B��G=����ϋ��\Av���`-2��L������[y~��o-:sl؍�>.#u /_��#�*���Y�{i�~�#��Iw(��f,��Æs�kA!�i�~/V���%]�H��Z�f��*~�.�m���7��j�X;�6�9
}�{_d�'�)�$H|e�q?�U��W���}��n[��j^7Q��j_Y5�S��N;˲�����Y];�|�2	C�%�7y�	Q3�<!���ET����0�2��[8��U�к��O�`2�d�\ޤ
f][���0&H�R�ޒI.�c<�V��C�m������ε�\1����"87|�C��	�˞�9"`H�Aγ�BҎ�@��5tj��F��璬���Q����4���Ώ|�H0e��C�� ���_k��S3^�}ut�.���-q��u�&���H��qƫ�����s�1�(j�H^�V��q�J^\�������P:�C��#��<�=}�`������o���3|�p�0���j0G��j�px$���"`Wٜ���>�)f�ǪS���ά�����	��v�&��x�"�҇ԑ����hy�����F�1��8�oq%�H�;�$��Q�N���8c�'耭e�ޥ���~�CY.�Mc�<���hc�P��]G-���Z��a�_�k�\�Z+���r9Y$����o@�$�골�c�K�P���P�h/�aG`{[�;y�0#�a����$� �i�rB��ꤌ����3���ܗ����3�b��r#�i�O/\���s���{��Qs]|�n@�vdނL��R�䗾>S��nl�N���(�}�+y�s�t3h�:�UU�Qz� &�B�-��Z8�!ݞ&?E��Vg�^�а��ܳm�v�q�d�C�S@$��%w�hU
����y��H���:�*b_Y��$�g�&Os��,����q���	ڇ�x��J�}�kw���[AB.��tއ�D�z�;���cI�K�/�2�f�)��4�.XȾ^��M���ڄ�HQ�����k_�g�����F��i~w�p�ɸޛ?�����I�ã�ByK��f#:�@�0�gS���4��	M�cb�	��3��7��G�	��}X���&��P����xQLl��=�6�
�ߣ�^3�Tk�j����P�h�v�J�P��u��isVw��Y�c�t�4�K���p �����ɍ���fg���D1���O�ن�mӪ�ū?`�p	(lAz�uH��3��������{�@�����P��1�d���PQV� 6F�
uX�HV�N`D�Efǹ%��tt�x)0WX&�x��j6���aW<d�����^�[�}P���\ҌS���ג�5a�Z&ɦ �f�D>�]�鼌z�A-A�x>�£MП��^A*iw���{d[�j!-qs�@��)w���G4m��W�%2=ē�L��@������k��� n�XaT
�W&��ܷ5e�D�|	E����g�=�فxY�D[�D���#�y��/tF|Z�+ҵd��
V!�P���'a
�=i�U��j|s��m�A"�~l"��]�S�س��:�Ƭ~�
��k�ש�s���T��@��V��Hf�K�b�)�[]z6�[��� H`D!*F
׃�`U*�(��/����I�G�y-��J:�;ܹ�]�@#Z<g����yU�h�^�E���%4�����̲����/�tm;+e=�t'�T&��j)���rX�,,h[���WxH�h)(A�&��~�q�ld���:�˾g�.i���X:�tn"jM��k�}�M�^.`>��\��O�KF��>�4�F����9�?��7����Y���\���~�Aܯ�#��EX,<u����U���v�Yq�/E����U������逽!���^�:�o��+s�ʰв��V��a�\�Djw��Ut�١K�� �(�2B|QSk0�@��[<�A�F