XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��SR,�I������%��ˮ��^Lov�X�Xy����E��q�f����0�ّ�]*����J�\W�a:vGar���T�b����R ����SKXg�	*)q���"a�m���\�4��ŕZ�L�"=�j\��yB��f��d�My�"�S_�~
��q`h/����k�+$p���
mi�W��'�	.�M���·$:T)Q��^�1�>"
�g�UV^Rtt��C��K��������m`Ľ��mF��ި-F����2󝯈�:za���`�F��o�h�fw��=�&�����ަ��R���@���L�9(���流U3�v?�������J�S>�����,�f�W,���ѹ:��������ڿFy�_Ƕ�Nր���r�V�I�Je���̼1�����ö���`����dLd���8e��W�x�0������������:��%��MҩCy!��L�F��؈W5\}a;&���a]����)�W.����*~JB^��aA(�e~��J��ѣG]��4�����VTSW����6</K����Yv�ϙ�@�Z��<���p�?������5�4�x��NX��B8�YD�YH	�1h�:wD��#u	w�5ȏe�m_�'����%����.s���
����p�C�uυ�qZa�W����c��������O�T�$�9k���g�xt��|G�N~�%g��$�ѷ�n̝��!|��u�P��R�ლ#�1VrNXfqky�I9Y�XlxVHYEB     e07     680�Qk �]f�#_��ݐ�XI�}s.�����clZ�s���:�s�x���T�>���'w��H�ɬK>�!�oN���'Ŗ�F`Y[X�� �#�)�m8��d���ߧ��Gx�#߁T,bخ��M��-VO�9�b؛'���"�V���u
H�H�(�/�r�/4�Y�����%����x�1���̧��2���v;�a^���Xsit�i�	<����R��ۄ�%�ǣ�b?ٲ��j���Hx�Wq�.��3��������-���] ��G�k�,���F�����}��Yঝk���z�J��`��o���PݿNF����P�D�#E�c	A�����؍�DS��?ˏ���,����' 6�z��nE�~j2�V7��E��x
n�A��(� 3��>s���t�1oE�D�8m8�����b/��_���*N�6n�|Ӈ��ܭ����*fw��jB�tHd� �3�!�����.�׭�v��z��"�BM�#�����:3ݹ֧����[� `�(���ʱ�-�xLڪ[["�� �t��&;v� C�V¾B�N��CSu%sOCcj�,��0r��?G�ͧ� ~鵑�h�q��Ȁ����Jc�!�7���Ѹ#����K�?|7�.T�*ޞs�!~�5�\�B��v�j����B�K�o#�bx\+o�w9_Λ����cBB�G�:�s��q�q�ժ�$(��۰e�s)�� �A��,m����9��H���K^P�� �L��6x���(o�C� �_m��a<��F�S��7���"�..�!�9�&>�"6�FW��^�HR�^XsRZ�s�qTkeF�_���j��-��}�')�$��1���r�`2W1�WΩ"�S��±u�P��c� f%6R_\@���Ғ��
��yu�����ЎY���	;|~c�<
��nP���.꺚� �962�<��utQK7[��,t�-&���Cގ���\n:��=���jA���l] ���xr	��a���]�t��+�=Z�)P:9Fҋ�Ge[�ؔ�&8�$=���b�0�%�pj��Q��a�4qݍf`�F�K7�<�pÀ	U���+�[�r��ɚ�yɕ�QF��59ʰ����d6��@�.b���շ�<���u��.�B��GR���ih���!��Vu���x('����w�[u�����E	kNtU���7�m��֙�D��v�ɾyG�Br;�\�;.+�Uc�^�Ĝ�z�uUG��H+�Z�Z񊪿H�� �/W�_�R����2я�i�#���=o���R�Ӫ���ĥ&Y�U���޿$�����q\�di���̝ <�`��W�R�R��YӀA�� �!�4*w�nA�;�h�ٲ\L�ԅ\,�3Q3��E�{�<i�m��z���_
����<�#��dCj[q�=L����YJ�I.89�/V8؛&E����XE�9Ҿ�ڎ�k,�M ���4��D�7���h�������Ӌ��c��JBGU'R�Ǝ\}��G��UOr_:+��]'���Z6F���#LdZl ߵ�7�j-|���2�!א
*�Xk�a�̴�N�
� �}��ey+h�[��ah�ӕ�#sA�0rk�<�T�9����^�