XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����4C(6����ԐB�d��d�Z�e69�����5_�KI>�7gb�tg�R�y��M^�i�h[fa7�RXI�<�E������J�{)W<�oo�L��y�}o��{���2���]�E� �/nb�D���jZߟ4%9�|�0�(����$s��ø��Ts�QtK	�ʲ��HǷl�J:�.쎻q��F���$�ۯU98{�$���j�"��0;�5�oV��Qi�J��;U/o��Q�ٌ��YH����
i?���dHΩs�/�H��Ќ�*�\K�,^�ǻˮ��Mv�r%�	.�V$Hj�62?�5�/r_�Š�R뻵��:泦"�`��с{���'��*TeL�=
/q߲,
�O�`���@
ȓĀ������?;j�l鉻��=В�d��)�%�l��4M\�������MQy�D���a &�F[���8��י��B8f6uu��Fi'�d&O�ݎ+��O�R��ŮhL)�?��$�#�T氝Ǎ�
C�����?���v1�%,^F�Q�H"���ݟx���h;��;&k�C��B8��c.�vF�	�p��e1��Yc�΁nx����H�UI��*h,A�W%?�u��]<r��FY�_xt��֬F�+_ͯc���� �����$T�/�4<�.I������#�8�P���o/��v�OO�~�.���K�t��p�u�>(�<P�ę\͒f;2Z'��Gd�x}(Lz�(؟b>��+c�_yS��b�a��T���kW%t��<(XlxVHYEB    4284    1110�w�ID蜫�����|�}$�֣�݊u�a(��*h�a��_�NHHҰδ�*���Y�Z9���v8�~AaD3f@�hJ�^1�p�N��.I�{-��t��y2sw3I��o��(�q���d+֨S{�OYL1��7��
���I�"د���7i.�$��Qʱ��1�X0���i4wt��G�#���1��W!��	��y�t̲��OA���3�nhZ�As�b{X�bj7z��ʪo�,+���'�>�^��Y�{�X$����l��J�ڊv}��KzQ*��q�[�W�BV}$d��6�g�L��ç�-����R����;��]�C�YJW#�,O��wS݂��O(e##b�r7e�d�I�?�%���;��XzN�+���A������u2kp�c��^� k��<ˬL��S8��gY��#Z.��DX�F6�)�k��zp�Dt�s�ަ�cfhWv��!5@>V�\�U��F]=���Աx�gF>07Ts��d�O����\��3��gH'���2�`ѹ!����0C|ڪW���c�)$h����q��Tav�'Q�����:@�7OG�H�C��q}��y���z��z3E��Ո� V�Z����4h4�$ ��R��d�G;�w�Ii!	�6>?��\ƿ����v	�(�^pd�L��x��Ҁ��&[�������-}��ʡv�X��tx,Y�*�Q�"����L,wX�rI�x1q^Ϳ��)~x��m/��$��iJƼ������؄X� ���s�T�`$J(�����8BJ��(�Bu|5"�a��s�b�I���#�c'��N��@o<ei%Ι�V�2e��|3���ر|5�����āx8F��U-°�{��jk�tt��]G�j�3;�j�ۦJv�H_�ԃ�NW�k'h�K�l��a<��N~>���t?����gi�>֕���>kU~|�fF�O��(p"�|�o������e)M���zPA~������*=�c�Uq20e�5r��.��rX�o�(w��A�<y6J9t(�Jb����Yh��|am��9��}�]VG��¾�س�[�ٛ�ڴ���>�o���\�L���������Kڅ���ȅ@7�?~�13��X%>�.0~�s]S���d����)�@�^e��W�JZ���BN������_��jΧ?�#݊aE�`�qrTo���P�W��so�7<8
����;�r�c&�yF[�$�8o
XEu�2�1xLjj5�MTӻԪ{�a���t�#r�AqР�w\`T9l�������smP�鸶�#��K��1��4<�eK�ݘ�1u�>�����ZkZ
��t���_�~7>�1�?n[� c���o��B������*�����ԟSO�f�xW�Oצ��~)�ƴ�kC�Fi�"�E7�:���P.d��^�I���{� X�Ef�h~��K�b��5]��'�o*&����C��ǻk�^��N�P[R��)��h3�pp��D�{�̐��f���;m�Jcް�М��������ݘ���� ��)7=���[��c�dS��O��dVT�4��L��S�9Δ
-�:���r�j��e��򋇷��Z�w/����A?��	ھF���8��HH�B�d[7k�p�MY�;��f�{'�,�8�ޙC��y�z{[�w@j���������{�X��v���6�Gۖ7R�e��P�H�&dw��\$5^�3�WS~g֚%WC���08C�����|YL�\�a�vh�� �e$�p1(~8=r���*Ӹ�-S'8zU�/(l7!+c�P�u���r�\�-����d��M���B���X���,�,ldS�s{��2�V9
�?�I^B���Z�n�|/�_(*yE�ȥ"�N�^<a�);�YI&hne��:? ���,�7F�W
�X�K�T!J����ڎj�֟�<~uQ��K���c \s�L|�R~H��eב`Bo	&��F�%���1{8�W3J������^g���t�\��@�h�f!61�ᤃo�������l�7�jp6�=���m~�������� ��z{Z%"����K���4+NCg�q�dI�Ph;=�	�D�+����,�=��m���]�d4��3�!098-�EI/�fIX��v��4�_b�c������Ag],���J��5��`�_�%$\{��O����=��)���_й��c)y��B6F0d�]$��a�x��-S�qUgk@|�t\vſ�2�b!C�
���E١�"�9��۴g����]L���������́2z�_� CT�,0,�OI�9y���;��X�Aev�Hb@�g��ɾ�yx���z �y������(<R����1�Q]�;~��Իp;�1�^�@��	�(�mg.��O��R��f���N�u]HLx��Gq�6*�|�/�<�T������[����a��W"`q9��a@�[n��<�n��ʽ���t�Wo�L��[EA���_��2f^��������ӕ���6A�_0�Q�W#hU��c��SO�r|H����\����Akk�-�'���>�`X�浓��P+<E���^"�x���dfJ���6�7���K����>k�7ͩ�w�6é�k�@�`C=���O��^b���Ll�{㇔�v�'��V����F����r�2#�<�4� �����&q�ϫ<2n�	��.V}���'1fxI��Y����;]}W�
}ac�ˏ�s��ҋ���S~f��	�G�t��4��I�<�[c�0$u#�O~����'��7��������8����cj50*�sO����B!n����Da=��v�wϋ?��*��sy9Q��?�^�ƿ�fG�د"3�Vkŉ.�^�W�Y�#V�|�U���\~��y|r�1s�U�k�o�*z����q^{���9��5؞��\ܓ�0S�o|�2�m�t��`r�������T7�ze�/u���G������r�UA��pp�K����:$�s�u3C��J���ˣ�f��j�/:Y�������S�Q��=�]&�^#�?	�3S��@4Ų����(o���p8_4�!�<m7�����A�(����
s���E�`�m��Cx�����7�Xb����Id��w��Ft�cl�u`�B��EB�L��f���*r�e���'Q��Oi��I�����J�m�O#jw��8���HB��3��A89����z��x�������i�|"O5I�"���������(hyb�ʮ.>C��[�R�<�����t��-��z�Bh��j72J�J�?�Q�K��;��@gJ�T� ���b䟳�� ֍�.Y�qr���UQ�h�';��64\�j�c��pOu�zeL%�3v;5���*pm��tBP���'{���:=�1I�O�Km+Ǭ� �Vp�	mo����/C�M��ށ=-����-��&��$2�W��Ob�+pv��k�[8�l��3#��\��7q�b2���ZV�K�ȧB7wO��d�j��c���5skH�1���݄w�	��ֻm�7W[�P�6s$��).�j�+�i۳�Dd�)M�p�^��Ā��"Ϡ��t���ʖy�fEp.1a��k��j.���e�[����G��GvY[�x!k8��l �9Du�����=/��ojźʩz;�GyP$�\1���#fK�A��)�}2���]�1�]o���ݣ�dQ�	���\0������ֳ4��
��������-�0 2f����[�=F�
ܞ��Of�����CSq�i�o�uc���긦�+{>�l��O	�n���d/����R��PB5n�=w���U'j��3�Bǚ�7�3a�u�:����������l�4�7����bqǅ�W;�,�oM��'�����P*�E�|��,�@A���irx|�����u�jU����?��}����j���?.}��������_�F���s�"�ա�U8��x��K)y�$�g �����HF��]�'�������؂��N��W=�M}�Zy_���=����ቲN�v �YP��,��2qa�*ۃ@JXr�O&�� ��192⎿� (��5�,���a�E��9�}ڐ�lOh9�wРD�5�h=ɚ��{����UGE�ls&���.��8�P����U��i��UjH�I��U��R���_� (ײ_����$��� �D;s�(��	��J�H�ޙ��E�ƌ��:qV�v�=DD�4�{���Wa,���wxrqN����nŒO"ƪ6��|}O�|`�u�U:yb��="�