XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����$�FRlYuu&����l��!�����E�NZb1�*��Z����v:}	���8l0iB�)��7�!�Tguy�6��&�Ê?´(L	GҨ��F���`�e�� �����
s��κ4{k�Jﾐ��\Mr5���~�:��V�x'���d�R����G���f���W����(^܄�3�����g�M�m��_�&���W!d��A�\�aG3ކ�|6��b= 1Ou�ǫ&μ%>Ն���p��#|��!%-����)rIʎ��Vo,洶�C ���Z�[G���W�OԈe0�L3�Z3�W>N�;��y��8?w�W��_PE^4L75,0c�n�?-�{MSk,�iٷG��5oֶ+�?��@��<T��z�(,��hG2���7A?�;�E��2G,u��	�qo�*f%3q�3��}�R�q^l>�&ё�q('�~:��2�y0�<giQA��Y�V�JT7j_�Qs��߆h˿v(9�U( s�Ҁ$�l�M���Z]N�3��i��,����#��!BO��s��	 e_}�kr!� ;�$)�_,�wb��W{��p�Z�����3��� ���t:�}�9��	_0��O�wyz�"�Y�h��l�.�K\˝^#���y�'��/���0x�u��W���� uZ/�ĵ�1��/9�[���+`��OEs�aI�{���F�rG�N{_@2���N��ݠR����}Eg)o��KE>{ݎ�5uu~�m~p�HC:~G*wx��D�XlxVHYEB    17d8     890�?�Y�RTD�Œ���^�Do_�Gq���&��*++X��_�DR���a��d��R2�-��eW{T�ۍL����~�����ĴD����Dp��̡2�tL�S_�B��fEH-(���CM��=[�!=*�*�˨M�U��w�:Ld�4et�V!���>���yCs�y%�)�O��,m�Ju��h��^y���ܳ��]� ��_�mQT��2�ټ�j?\dǨ,��'˄�U�@�

�n%d�������������f�����m�U/���
����8�L5��@��qj%Mԑ%
q�}�(����I�#��-�'�N�`��-���Q���Z�n|8��uV�v|kwW�q�����<.���i��Q��t���|�h��ڔ���
]���yŮ@���Et��z��c��	(���/�G=j�l���dH��-U��2��UF�*�<QձZh���-F�li��?w��v2{����R�F��[5ۣ#���ܙ��U�:_��&Cr���U{�rhR���U��ף]�=g���n1�rLrUjq�]�M:�]'�/*��:`����ͥ����"�e?*1nkE��ݫ��c\I�m`�����Ƽf�J��4���ю��������rA�[޻���� &:Rl��+i�"�����DI䢠_�[���R���&��\�J_1��
b�>~`����S�WbiF��8
]�j1�L#ڮZ#)I�0k�X�� TY��so�q&O �ɹJQ��i�+�Z��o/�XM|�7�(�%h*y����t6r}I�Y:��+��V�82Y�d)רӀy2c_|��,a�Ѳv�}p�9�i}~��Mݹ{�bZ�d��/�5Rn��Z��LG��8�fD��ϲa�j�%Mq�6C�P�����!)�J��s4�������@�=��~���m��	;�"�Q1V^v@��s�=���O4ap���K����9͵��Hy^�7��n6��bx7�x %��AA�� �cBWDUl?}���jԢK4%1�@�e�|1�����@A��/8��l_�U5����T�t��;�W��gհw��V�ix	����K��ܧ�s��}��ub����}�=���80"�����R�uD��Y�_�6/���/f�A�3��\[��߆��̧|үHQe�e'1�x���a�(�l�t+c�_:�����F��HZ#B!��T#��L����R/�@����)��.�Q;��~X��?m7���)������_C�����ː�
��ش;�O`�dW�M��n߰�
����0r���&Ό̉��`i���<%,]ט\R�p��	q�/�?HLz*�5Y>��z����\���A2�Qٯ����;��T����zO���l�E��S^�f4k%u4��)sqd�N���5�(�@���7찰ډ��>,�k��D�cc�;]�V��ym�}��i��>�E=M�-to��+nb�FI����)^U����̟���P�	��/WP��i2v_�<�ܨ������[B���:��O_����6{�6�BI4�D4�>h �e��G����hd���T���؏�T�H�� �V�3$X�p�����>��^��H�k�����^�	l��i�@�ϡ͎�ߋ����u� U��@n�1���is����2b3�̺�A��!��؅XN�bU������
�������M4.^���/�;��my�C����G8���X��ϳI�{D#F��gŜ�ɢ������<EG����	����� ���d,�y����^����{`�'��:�#D}�������^l1��p[�Sd�x����,s�iH�N�cV�¢�|W�L#�! DX�l�a��|b��J���/:?��t�$�f��gTN<L\�&˅���P^n}jN,	��n��N����,E���U�����y���!�#�5e�*����5I@���V1����c�Y�Ϗs+�dxJN��_B��z�A�o>�F�����Ϭ$oC׃�k�<6��\�6��
��@%f�'MW$q�P�r����٣��l\�a�$�%�#J$D�S荞���/�x��x�+O���Nm*ɪ�~zq�^�?'ݐ�O6)ѻ�~���Niv�e��y
�˸ G�� �g#�#Nk\;