XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���P2s����π�����z�9��p�����G���I���18��O��ğ� Q\���9���sC|]��_�Gh:e��T6�h,��mÉ�d��0V��ĉ���AH{��Ԅ�-_�  �����u���yea6ЇU�'���W������0����Cf���t��5ܸn��3�W
�2�;�ͫ����UGo�}v5XF9�0C$d��7���1e��kU��7'}�xs�x�U�qh�q�;j��ݪ�J�$O��{��O Z$ Z	P����R$6�`ᑢ�W���s;��6@�����z�g;Ju}f�XӎGt�,�./��Id-�Z�?�۔�]*�Pjx����:���Ƨ��lФ�����v�k��Ӳ�-y���_68�4R�W���G�k���o�4	tDwW6��d1��|�Ȓc��욣��!p�H���6���`X���+�i�R?r����ʝ������k���IV�m���}pur� ��]����|u.d��lc^�#ޡu_��b��!�?�3(P��Î�ԣ�o�Y�	�\H,پ�8|�\�$�o>���K�C�V��i��4��6���Ƀ�+QxD�I��J�#�Ft�i��۶Ѡ�v���)���A�29P�4��,z�֤'�$�Rc�cC����6�D���	��ll�����)fEgth�)Q�:p���a#ՠI�[������f��h�ȹXխH��!�d2�1( �,'i�N�hXlxVHYEB    5d29    1390��c� �Y�Jyܣh��k��QF'���n��]E_��C��I�;XWW%@B
Gg�%�k�9-_*�6�:��O�� 8�����?.�Gs�N��+:����p���U���������\gnR[Xq�/�r�HeC�t��ce�n��FˠƔ�ًB��a�ϒ�y�.;{ta۾�dH���A�׀��.���Z��t=�Ny���>>�t<*�*+N�����gg�	�z��0�?$�Ll$͎z�oն�zЕoU��݃*���>|�t�8r	Nѻ<�S4#�#���k��*[�<��{�q�]xN)�|�%��	O���r�f��-�����wrc��~�^�6>����.��s=���cHfr"���F�� ��'��"B<��I���a��t4�qaTv���T�D��@�M>�~/S ��A"����������	cmw1ק����{yL �4^X6�	��4ߪ����`@&�\�7�눓���������RA$i���R����#*+����k�~-P!v�*BLr�u �,�U	32�%�G����w�*8��#sE�����ل!���p��^��~�\�h����c����{ƴ.��SM�9��Ȏo��W���9�ѐ�ꧬ(b�w!4�� ]�cH�~�GAW ��za�e�5�_{�6]-ӀZ��]���a�&���f���Fֺ&�ސ4e?�fA���wE�p����^،,�� ��Ń�h=�� y��=T�6�6R�1o�c��,� }k%d�	�~�kV^��K�1o��cՁ��?�)w�puﰹ�P��I����H#@�9	�*��Wf�x���a�_��i��8�Q�@��W��3�I�N{��@x�T���cJ�����"V$��y�����JQ2$KN�*�ao�4���8��{a�"uG0Ř];5��a��h����c=ܬ�,��l.p��O6��U��@;A��+CCǻm(���{F]R6��!�^����B��9�/k�=~�k�&�>���B����G�� �(�h�!l|�����������25T�%9��`�m�ռ��Pˎ�=4qtፓ��%��yN�N~Є����iQ�S�������5@Կ�������s�`�<��tE��B������ѳ��A��G��=�*�U��]��*���͢&�=U�ѧ)FX���J��Kl-��e/y�����S&��:�b,��_�kFn��Ȟ9R%�/,������=��Jn,w�$�GNs?By$?�ϒ�8�����φ����{a�@f�%��#�h��k?���-������u��H��ef*/������x ��"�\:����迶\FÂ&)����c�2�wS�w�i봄�2��A�y�^S���G�\8H� ��3xdC��Ú�lUZ���W'�;�w�u���dŐ]R_�U�ܢR�]AI?j�m��[=�T�����R_u���?�D�����r��A
�������]��	o��ňZ�:��	��O7'�܂�2!N����K_gb�g�=�|���.?b��^�o`T���t�h&b���yrBu�����kgYn��%u��ǵ�~�X.f��
�i8�j�����h�V�	:��Z�!�\��r���)��WCɢ��vت��AV�*��l(��C,���-}��p5�~��j?4]gۦܧ2�S-� ^M4�Â��w�V�X�S/#�,����g���� ��S�	F��J����C��D�e(M�8��_W�����%)�K���3ს>�}	�&Hk�]B1w�Æ��[H
��[���!�]�{�)�^�d+0���	��U/f��e�P�v���M�U��9�|w빩�����s���h����s:ל�?L�x)��:�x�x���8�ag����N��+������QQK>�r�����u$�I�-I]�|�$ǀr�����2:2�u�?=\yg�I��[���N�s���)�� ^:g#]������`�?y�#;VE��B��,���(�G�N"6��8�:p_l��p�^���T؝&-����@&�$I��[̺b�0������"��4V���W�U��tT�	�p����l�^K�� .��|��l�ʹȼ�p��I{��eI��7����~g*�N�r�&)�FLd���?���f����=h����zW�)�����c�C�p� Q��ms�aq�O����sQ{6!�����m`��o%��K�&�^�/-�u2���v���O�[�5@Ŗ��Ñ���C�u�ЊQs�����>���Y`+�G���V�'�Ֆe�,ԏl���_��)��v���e�VB�:/?H䩹4���%?�(�5���;TP�� Q�g�6����dk6��SM�p16Ja�$�I�wWgpB�0����-{��������/:���l[������@C�ꥬM��$�ӳ;�Y��H����$̢�!W�6:�WL�P�ӓQFy6��ХW���d?K��w�=�P�RPK��͟��W�B%]|�;����tRa�A�R���"_\g7�E��~���pG6Rѹ�鄁 pY�![�r��V�]�A�/����iQ�i>p�~�G�c��������U_��,�K�bK���4�q��n�e�
cț�-C��;r�4���k>�/S:�ϛn����'���� :I#/҄V7�wgը��Ӹ3�Y��ғ�M��#SM����"]RcO$��@��?�x_�L�{�O�Z_I⇍w��5`�p_�F%���ɐ��|H&���A�`L�#5/�P���5�F����p.Jn���N����2� i��_��.����A`�s��јٺv�Ku�~�g�r�8�J�ǣ����2��mG7�g��b���u�Ƙ�!Ǒ_�b��a)����Uǹ��O����ҧv�t~M	<^��K�����<x������ A����a�#�P� �"�]���`}⥻��/������A�=+�o7?�7�F�J�$�*ޕ4ɝû����.K`*�0�װ�tw~�mZ��W�����U�hEzV�����
�|}Og�H���0{J�Cb�+1��4�Y�>\y+�:�Koi��N�_Q��Fv"=�_�q$�Z�"��*����V����㔮\�bV�6"����Vy���w��Ƀ�����\��Df+M0F�?�k�Q{'���71�Ň�BD6�Ɋ�u���7�7��?Ϩ18q�uӰ1Qm7���������0he��S-7�5�P�N���I�+U 2�n���u�����CO��~�T��V��R����I��݋+�I�N�^m�z��6��b�����/��T|��z��n%�0�:������<��a������EVy1 �3G�;I�ge,�}*����	�aڗ�TN	MyH�H��T�@���=y&sώ����2|?�CY�� 0~��0�Q,����?m�
�)���-��liV�L'�$��(�;��2�m�.���;��9��}DG����L=��b�^�f�d�)Uf.�n����/ɭ�^��aKٕx�~yc���8��α�Ũ�iY�Ռ�TgIK�	�Hۺŧ�O�c���I!ah�P]nhr�sD�m5(��og�pFc��1/��@�5p����Z	
ړ��NY�� 7&'|��4�Q�:X�X��@	1�>C�.yGl��Z�J����eÂ(�n J��`�ـ*d�h����y�"�}a��� 1�3t0F6�~e��NL<[��9n���<#��	��������C2�,�W���M]%z�V���iCGd��a`���ͩ����&഻�s�V%�@�$��@���&��wU1E�jH�r�74���L F��J���7�mB2��� ގ�����v9����Ԉ���� މ�A��9�ؖ��v�N:�6l2�<#"��D���YIS�&�Յ�,���;���l���7�۶���g�����xꠎ�ۚW�\_�}XNn%�^�y�fv���R'�B_=�E��T�&Pq5P:�V����t��H���87(	�gl�[��Na��Ò��:f�7?�$��1�*�o�cݝ/��x��\�*�л�oJ����k����y����Q�����b{�f<|�����9t�Ox�#���
9|D�����4�=6�r.�W4�9)���[5KM����6t֎�Q��r)���JW6�V���h�h+�)���NE��x�q�j^��mk�	U�O"�������g%�v�������� �=u���*����iof��Hv��t�B�t1�j�v�sz���".�D��}@C�vv9���L[�˱U�0P)�G&4X��]������ukZ�h�mG�=�>3�5�J�fK�zc̹$�$��oM+�v�J��O|;W-��3��C�_B;�Q߲A�L�6��%Z��1�����a(i�� ~�ЉqCF�;9�/\�2j�0�PԻ�����l���ϨGu�"�ƣ#7�X���MJ�G��Vܚc>ꩭl�\W�(�BZU)�&�ϔzq}�N��sS*�uHڽ��N��d^i�¸�Knz��@YD"��/jk��~G"���sz��i��!�+գ��%���0�Er_ҜB,At;�z<�*jG�.�5����Znޟ��`*迷�&9S�dR{@A)����5oX�d�v�O�ix��tD!�'(Iu��#���OA
!]_�0Vx��g�7��YjV� ���a��$PL�q�H���w�|J7 6{ov��$��7���D�P�m6�����L?�7#�����_.�:T��������kxX�7��_'7���Šo�B("!2�2�VY����dGo���P���o���M�r�@�S<�����ǽ��FV�g�m���#���&�EH�<ť)(u=o��E2h+���Vl�.��+`�=��v��