XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����҃���9^GB��l:��L�/@�xF�#�]Do����,�py�"@Z=]S=�U� a:r =Y����~^�K�۱��F�#"+ǦlY����Y���ԧQbEW��4_��*E�c�6QH�s���[��8{��S6��0:>�i�aUkv;� ��m��+��M c�tm��-3@]��³YiGmMh�)𼵟:����}�uǵ�n�|b�x��vv�I�Uh$o�$�b�fh$�\Z��e|��r#�%�`f-}��( ���N����G�%Ӵ<��n��}����e��j?Ts��U�DKq˯rJ�T\(\�P��Ku�p� p*�㿏ۧ�T���(M�p^��e�Ӂh)��A�6A���Y���;�f��N�j���[�?ĒT<�R����%�ݬ�0=�jM�c���`d�v0Nγ����<-����Ҍ�L�S��gq4����/$F+<���h�4*�~ɽ�}�31LN%�'�2Cf��Qѹ���O��}����4%��RT����T��n������LB�x�뱬�� ��,��d�Z�3kt��ϼ-c��F�Y�{wx
	[�3�z�KFp���}�=K�e��d9I.h�7���7�y��U���=��FK#F� 0g<�L~�������PhM9�Q�k�����
 �����.����?bP"8��T �w`�A�v��+��`NZ��������?l��+	����{����g���ɍ�܇��v� '㭷$v��܍>�咮XlxVHYEB    1959     920Y��a�F�Ӳu��3�?�)����.j�z�fE�>�ӏ"��Y=�5ԋ���#>�x�����r�ޱ�"�8T���1����D���4��̰FNb�~[���x��+��T�n����세�Z4(��K�ȍ�������^��i��L*h��*�������qR#O"=��U.����W@�c_!����խ��[ -����qBj��w�Z>���P��e_ (���l�Y�}��t{�Ӽ[��H�ꚪ!�:g��Q��(8=��цn��X<T��,�,v�R��21��t+��!�9���2�w������F$׆>����rAP��<�xa�ϙ�������E�hڒS�/ZsB��Z��w~��X�i%��x���/��~*��1�b��H���yp]���HtEY�j�@+'qE��w�k<��-��t�bW���2F���}@��g�n���H�21�ظhv�P���?��j�L(�����զ1l�/�J3[��Q��@�V��s�V�WNLq�V������Q�,5����REc_ԇ�u�����B���"�'������UnG5��\R��+�O���\~�[6^nc;U1�� ��TJN/]'�6���ch��0����bT�����y��ΧT��H;�·����i��4����a`n����c��vz��C̶5�j����t�˺����R� ˯��q2	�F�cP휛���^lPV7w��c�`ѣ�
Uա���d��*�����dV�> �l=ܓ ���7~�wEG^�c��Y��N���x DG����tfp�Ms���]#����φ�-rV%���w-�B��BP��my�8���%����8�!��5w/���%m��S��Ԩ��Q��w���l؋�nW$���=��ϙ�OK�g������E���1�g�9��ﮣ��v�$s1dfV�ר�2�x�h'`��tB@��.y�e2t�y���l!��f4Rm��+��Y޹�,A�����9�&��m��E����{��U�o�B��&?���g<�w��wz ���:lm���ea�r ������M��DÂ��9[�U���?�á�Ǎ��}w�,��#�J��W��-;9��6���g��i��3���O�kp�+�
b#��I��(�@I˵�g�~§�W=Y�$u�����k�ճS��� �YF;O�<�z�ex���i���z6��hA`y Wgu`��[���?u����˦Ec�9����UE�o��v�Oj�^�$'�T��m�*β����?�`�
����n��y`���]��!r
�N9��m���Iw�kv�,Hd�_����mO��\�����m�St	�i����Xލ�G�Mk4�������,9������)&�6��x?��<d��R=J�dYF����Uql�'H�]�0�.�RΠO&���3�I�J;U�Rrhف��U5E.���֪lT�] 6�'�*��Go�X�\��v������N5\�'0�1�Z1ѯ�ܲ��Ը���Z��-0����!�6t+�(8��X�S�0��+	����lWH��َ��]G������$����Z��+k�9��8�s ��FY�ȑ7�T���s{3Z��rI,��`d���迅ّu�sƄj�>�@˸K�kU���z��I�BE��m)����R��l� %�x�F�-����:�lK5}�K��`5qX�~y����Κ��X��_����8Pj��hVoy��F7v��Q'FBK3.��3_�C`jŨO9U�	ʕ$��/H�x��->h�ba���fo�u��	�&Lv!���J��e�C/�]~����`w m���,2�2�I�Htlℕ���q��P'$Q�eA���P�}َ�xe�2c$d �N��p��n8���,cQ(Z|��a��-��U9��w�%�x	���������*2_���+.��T��_�mjy95a�h,�)�� �ph��z�@��ФGp�ɋS�=��G��̇(}FV�n��!ꭉ��0�yn�g�D�D���k�Wpނ8n�35l3�OX_��A�d�V���_5q�u�+J���]�X��N����sI0�s��m�N���0�ő �y�Jg=��]���6e�ڔ~̏�������S���RM.���9�$"�@M��h��!BD�Ŭ2酝gse��E,�(cX|��_��Y	�'���:)�4ڒ���ܗ:⸈e�	c�es_� �њ���6XƏZ�O_b������Fi�%�|~ٲ��ډ��z�D}fcKW0+F�9�۳�*��.�ea��5