XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���}a�[DZ;����>v�tR��#�����?�����3$Pƛ:n&�M�����A��H�;F�(�v"��1"Ck]:�9�6n/Yd�k�?���۪�a)�|-��~�R���b^���A\�[�R�9��<T�4ݲ(�%�����4%ٶק܎��g7��({��g�O�K��h����'�8"˵oh�Ҕm� ����:���R���82�Ȏ6��f�ª}��z[_a����U�b֮p�k�7��T7��2gK�G$B�A�o�cXBixQ�\G�z���"�䟄:������8v�֑A�ID�y�TH��8�쎇1Bw�ݥ����WJ�4���^�n2�,�m��F��L�S
�$�>Pшz�_I,�3r�P�D�����=^�@Lm�
D+m�tL�^�ע��l$�+�q�ê���ܐ�|kys��'*����߸�_��F�03��7�۶;r+ �*��7��u_�и�?����]N(͚k�?�XFli
'�mOx�ɉ���Kp�9 ��&�n�j�.�Z�
Ɵ�[��$ӄ��@�#���"�J�b��y��Fe$\Y9����7����Gdx���T��`8�J�4��[�j�,8 ?se.�у��}�g���"X��&J}��䆺 �a�;`�e]�V~x�����XUƾ�Yfn��ł���.�ֿ��Ë�����$w�?!�C���Yrܓ��!��]��s��v'��b�� �RĠ�F���aE(&z�e�C�
�TF�TI�!r	oU�^XlxVHYEB    17b2     880�UCKX?E�x���k�d��*i&�X�A|�����p%����d�fۧ����u�Aq�-_�K�D��*x<���ԐB{�9Q9q\�/����[���	�)\#��<W��[���^�Ƭ�J����h����BE���@���7��/�+/�8���=j�a,$��c���ϲ1�;��&�g�����"N.u�ɺG�<���UT���+�D"�E��xmn� ֆT�?)��ԝTs�M�H��l���֮P2Ur���we7DxFB�wJ�Z[��!��#�=��R�N]�f\�u��	9Ҧ柤�'�!A�WsEeڪ�Jh��c��(_�{�οr@�|B.������!�Ut>��.�K��_an��]V6Z�I�
�b.��	<y��j��N̑W��Q�N�j����/�k�#�����`P�8x�"W�>*�}�8.����4�d�+H�⯉$���c����$0)>!�� ��"��q���S�#�!V�(�B��VVҠ��`��}��m/�]��x_l.�I�Ps�x �4���UȜ:n'�-�7��󭡥��#F��IL_E�xm9On�,qV�^�g�n�Y�\�nV3��1��X�n�7!�u)�����؅�@�*]�Dc��kH��bݏ>B��������U4�y ����Jh���U�����5��>���B%�����/t��Ϊk~�p�Ǥ�Г��H�S��,�ƹ�G�V2a������d��ڳ~�6Է6,M}�J�D'b�U��a�$z��z凲c�\A�3��Q� �Yb)o5kP%������$�f��+�A�kj�jw���֍��G\X�3�I�ӽ"h#�ܬR������z����9�!����Nϰ�q�~��K���Q$���%�Z� ����R�%r�L�����"cz֝OK�ы �1~�ɾP�1���L�
<�|�cT�+�`�c�0�~��	
��2��a+��y)՛� L���dy�߃!�N�o��E%.*��Q�?�rhd���8<���M	�3�C+�Rp�o{'j���_R%��p ��;7^�^�z�u��a�Q��{�Hޜ�yͶ��y����o�%6�djԧ��}���5���.��֯��I<�T�<�5�MzpN� k��������{X�`�o� ~s���̥�μ?�3��+������x~��v��e��P��1��MJ��j���m'e0"�ͣ�ڋe�l�R�X����;��e�e;Kq��R.����C)*�q��p�&��	A�%�=�Hb��׾xRLb���xC.�����Q��-3[�}��9�V���O�~P/6a[��g���������h�ڰ)SlRM��x�?շj�K�al1�!���Z�AIe63,����FV%<J��q�r�GD!"-fLD�S%ɣu��mA�j@t�8�=m�g8�o�.��]���D6o<y��y�礚�4
�pT	
iD�����o
F�>���e�)[뵸�J�g3Q� ��2R(���J��Q�Ci@�a��󵿋$uc�nYP��X�(S��W`JC���(��J!�C���b��^h`��Y��ٓo{2�y���G��
��[�Fd٪~�����w�b�X^	�+�����%���=B���Yc����	*��;m������)qF�@�5zq�`��SZ���<Anۊ����S��E;0SşbÓ����1��B�Ëp��v3et~�����|�IE���t�\��)|�40|I��]����P�&���6}(W�'¼�ll�BWkz�%��q����
�Z�*ڕ��.H
����R}Ԋ��ř�"��F0iJ������H�g��&q<��9�V�vEg�;��g�u��X�M������\1���gf��Ū��a�C�����J�{��x��+�bm䧃
�+�f��r���G�:H!f��/h(����Khs�L��� �;����oԖj�����"� ������(T�B�p�<��
���/Jdh����c����#,��%�G[������	d�r{�^�K��3˺U��αD(� ���gm�T�fy���.Ә�Q�J]��4A���
W7��6G�ڗ���Н���F�m9��W��u�񴾥�