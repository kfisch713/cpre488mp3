XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���K?@��X�m� 7���JvoQs�][��[L1���j?��o�� �s|�H���p�*�wW!l��b�������s�c��#|z�"����j4ZP�A�𜖢f��1�F�	�|x�v������r+��i�f�(�X�uu֘�� �=`tL�*��O�9E��;f^Ň�?����LA�Ë���qca7���$wO�(B�E!�*z5�s��6�YQ3��dddr	��cx2��$h���'�jl(��6�i�J^�	Ω�d���O`>A����ئ�{
!m!59I����H��z:j���v��M-�h��ɹ)�,xK�1�j��+� ��'��
D�������.ȩwZ�
�-5<����f���A�1`U��U�k[�S�ʥ����r���%�Sg{�O� ��^`tԘh��ʝ�#�5[�����X�Lj��]�k8�0�K�#��QO����v~����q\q�n�>S��L�%x0��C���u�y^W��{w��X�&�e�f��'�j�`��G�Kw��|!���S?gRS�@�JgWՊ9%������D������Pl�&��'|h�!�u��j�n=���~8i���8�L+?�Dx���+Ƅ���	�������xq�D��L���/��G��7���u�i�9d��x�x!�!Y��	c�00�7����(��<m֮$��������_��Z���m�K+~�G�Z���k"ܛ{3���t�� �t�[�T��7�XlxVHYEB    1959     920"k�b��΄�Ȟ��+���$Ȗ[��W	V��xhN�W@$��ş�O�h���&�Q3���0�zml�lw��ٱ�E�nW�u�K�G��.�읺G1o�N�
�e���u�*vebc��Ͻ�u�E�nşV�{��Y��'x�aq���6�t`:"�R3�N˗�/��#���ɖ\i���CH�*�%�5aa�{�;���� k.L��ϫ�g�|v���&�6ۖ��X�rg�L���j��:�z��؇D]�F���(އ#��ݞ/;�����\Ի�*Ӿ��@�4�7�5�K�#��!%�<7
��q"���i���T^t�T��h�4��w�K���*�$��1
�$�/<����]�����4{X�6�EvL�{0�EIL��3٠92s1�_I��~�Nm�b�;�!�+�Ĉ�5�?�H;XW�)�-��=9 ������E�y��ZB�q}H/7������P]�r��}m��/��hA,�ƌ���k^��Q������E6��&��j��3ަ���5.aj�&z����C0���w���65 y��$�~DR1���h΅*���)LI�b	'�_��J�m�!z2f\�k,.R�e���j	)�[��)=����-��[W�Xcz0�ֵ@�i�!U�u@$UKF ~�Fe��+1�dH�$%}/
�bI9}}QL�j��1@m�L�EG���,xeư@l��@���,��u{���@Rz����z��3t�����o�.r$��6'Q �F̗]�PcM� �Ҳ��m]�8���j9^X���x�1'��c��q_���w�P�z"��RX�p����l�A�$����?È|��1Li������t)5Y�.ֲ��0��Q��z�'��;J=jHQB�r�ӂ#��.���խ�1l�\�Ȇ���7>�`ѡnT��i���������H@���ȟ�ku��%��-Lz_���G����L��0�W��O�5.�T�K� �Pڡh/�è�|!�r�EՀ���'d(V�GR����:zīY8�	3�.�]��5?�;�Z�u����-�����D��:_.��}�n�\�S|
͊��:�`����^nA��P�u:&R����esexz���g�#���E�b�MZ&W�����N)7���E �<@U<Z���!$Y�3�'�%��x$�d5z(ǧ0>(�=�Gy\�;xKk������RJTx��|ك�r��LvTHh�2� ���t��>�����������ڮU�ddo�Ҝ�+�<Z���`���u!�����rTQEA�v`���}�����`�6����x=�39��ej��E�l�M�R�q.�;ϵ	�~�(	zjZ���%1ׇƛ�]��֗��$b���6�Ek F�b�V��G\�yܬ��.l�	����w-(ߤ_\��*����ynI���{V�#���DD�>�H)'U\��� 7��㲕v9XI�1����M��!ċ�m�&�X�L_��k;i��
l�ҹ�w�SƅհB�q�,��{�-o*5����[���DχV�3�u�?��n!�=�ϲ��~�kxcX��za^�$e�zX@t��p���d6�$���.�9D��˱b��P���b���%alӡM��_\Q.���)����K#4�I��qӅeI��AR���Ą���W���a�{�6�4Q	Ц��4��UՑ�����%��B������h�,�Y��K��ͼ���ؕ3l�EJ�����
��,k &�':��WCs{q�|���Hz�?�8�y)Ӗ�����np��_j�Q��b$'���;i	.�/*WD)�P,��
�V�\ot����h{���6<�IP��qm�&�Q����$��%P�e`4���;f��1&=��:�?���ؗy6�a3²dg�`�$��?��z�z�ϯ�~�T��x�Y��4�Sqo}�v�-tt.�b���d^{v����0 ���U��CZ�~�Q�����]k��M����W2��8���m; �P�)�H(@���@v�fB��[���*�ኁ��z�ӣ�F�V� y䕟ۣr�k��)}Uaz�:F��'P?z��sgX$����)r�X�ʁ6��m&�2��p�|�T `)��Z |�d\�w�ܛw��d]�z� ��[q�9^��a7*���VI7���$X{�$��''�����с��#И2]iqL���~5��0��ؤ-�?�*/�F�[�n	�dq���*al�HU9�袎p�~���Z��*�$���IM��6��˲�X(�q]�����"�������bĕ�0y��C��̈́�