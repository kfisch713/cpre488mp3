XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���Zh����$�tne�=�`�}BVB@	O�e�'EH$�G�0)���j������U��m�N��T���%D�0Ni�ۍfؔ9��@�fQ�(�YNͲ��3���u�6�-jV8#��D���,<��X)�We�����]i�ju\7I4�p+������ɍӦG�F#����!���.פ~H"��ˮ��%�������"�Z���B��)6;C}rŶ�����ᴬp0�����J�q+Dwrk1���'[��M@���1���|p�nH~D(��Y�q�g!;v̉�M
��tO�1�����r�����(s;Cz�&K˫E��l[,�|G��"�ˁ(�T�֨��u���� �+	���6R\���O�1����	"w������#�jܖ���4E�b��g����n�0�C}�B#��5	�b;m��k�H
u3��� DDԗ�Jq�ɲʁ�|�?J1��`XH&��L��<x�����-"+(��=͏�bau�[�/�W���oϴ�ql��;�x���%�u) ���,\�&�/K�:�����2怉�ᤰ_�Մj�+KY��us�;���G��o��s�تEKm��U7f��o�dE�����q%+�f����T*��}���K䆪K�=&�S�iWB�W�a�T7������aTf����mi��T�^��Xl|qx�I&?b��X�j��ǋ��ۑ�8*��p|��`�>�ѝ�7#o����J�Ɲ��4G���ƣ�'S�Ų\ԁk�	@�y�MWXlxVHYEB    5866    1100�(N�JM"��
�2�ADpǡ]2XW|t��_u��R�y���
�h>�[�gz��"��Ћ
E���x�q\va��?�u�'�{9�n#]��*W�K�E��~D!�R�S�Eq|2�j���R�:z[.X[���uCK��n�+��3L���1�^��'�R�@Zar�h�UFp�o��+��ʜ��#��ߨʑ�`����REZo亩/�j*�efNx�x�9�_��A]���O�2x�f����mrm��_�7��di������8��J[D��[�ِ�C\�:�z+)�:����S�����g?�(���M�>I�{uy�I(F��h��Ɗ�0��mM*N�:EŴ��Q� ���}L	����<�n����}D�n>y�޳��⨦|�26s>|��n����:���K��+yZ8�a�2I 72�t���a��a���5�����sj�75�A
�Ѫ�4��t�W/܎�|[�QWJ$�kG�B�U�(@�j��u��$^���ˮ��j��0�kVfa�5�����0}�G9�uI.��q�d����i��"�`�$� ̎aQ�6��<�6�0O
��7��KM���7�Ԯ黣�s�$��!�8�,bN_F{�_�t[�5�M#���4{�Ҹ�Zm�$B��my7�ۤ�9��� u�o��1ZБ�<�qA�������y�ܖ.!���I�>���	�O�W�*�4�c>�����Ü*�3x�$|�`M��\���P�}��)�g�.HK5�c�Ώ#�? $ʪL\Q��2������40mf�N@�׃�l�����ٺ\$t�$�BPI$.x�H���)�f���p��vY�O3�=f:ѯ'�$��[Z^+�~Q��-;���ʅ��'.�:�8u�j��"��I�d����aL�TS:
�0/�<�4,͂��T�_�5�`mݓb�CƠ�|��c�HC@�	P����1`e��,]�B��A��AR4��!/��o}��/$ߖ��@VBṤ��POpAD�����*\7vF�T�?�E[�ؖ2����h��0V&h��i�}4ITB`Kt��=$���N�]���EJ��հYTdO�3O��N}����5�4�]�5�.�o��ڮ�����8���m�{�oH��X���eE~�.٫�'�e�;�v���w�Vk�gp��z�C�������3������*�l��Mq)�-|m�3�?�,N~�;���;e"5R~%|��R�Z�o��4�;.���eL���"�2�����7x���^�� x�M�ɫB�e�,I��;1� x�,���C�:�7E��m�R��lQ�\��S>幆��g*�����e�t�o�p��i��Q�`�N�:�c��E]������0>��T��a ��v������ ��$&�_ d6v��8~o�`���M��oP^�g�Y�a�2{�<�-J,d��2E4��r`�������h��IFZǍ�ҨϾ���J��>P7n��[ZQ"DW���Q������w�e�i0̘ψ�Pb;;�0����$��(7��CB������3�5%���"RMگ�+R�t~1�g,��>�<#�;�ئ��:�mċ`�4��j�DD�BC[�JT�Pe�3A@P�=W��N��dt[L��#G��e;R�*F%���T �Y��Pv�X�z�FJ�/;�1�pB��dD���� L�f���ot���\�c��2�����t���w"�J���ǁ)<��z�+�y� ��gw��8����"���;�<jd�UurZO�8¥6
9����y��l�
�'��ˋ[G�q |fE�O<���?���q츈��`��PJ���K[γahԼC�v�}TNͮXZ�L0F��j�s	@�91�b�*�f	�E�Gq��=��9T9�ȟ\�n�L_"�5o�t�^�������A&���e��E!�Vbgl�wD1e���Aؘ���+�T��F�v-x���~�PJ�@z����)C�]BÀw��7Iٲ�r�7S �T��$�3t3�͗]̇o��U�jJ��ED�x��-{��V�]��~i���~��$Iv��y.�i�ߑ^=ڤ8���0�Tɽ;]�!L��܂%��T�߶���A�?p��թ�?.S�:n*� Ӭ�#���2�3���<ve�,���t��m۫�0�ƾ��q6rI��HVv�h��z�o.2�4��l��F%!�NM�,~���	�!��� ��r��֯E�f\�����7}\�6̽b�e���Z8�1M�_�:Ӗ����࿷`�k�8ǆȤ�AN5��b�@�z�����t��?��Z��h{w�ݰ�	=`l�A�~ގN#;������8�0`a�}KW��|�ŢJ�������8},�8-��z��~�9`�Y�D�	' �+�~�E��׎�r$y���hB�l�=�t��G��ͳ�0nt��l��mP$�{��r�<�.�#1A6��C��O��T#"��4U�ȡ�t�lK,�w��<Ƒ���[�Yl�!���6��!�",L㩖Ճ:]�<d���u�ӫz5����e����� �#�S� �1�.��p��Z�������vfY,�N$ER�3��	�-��J���I}�4��ю��������`2�'n��30 �����uy�i�#�|4�chV$h����+�r�l�����l�nb��R"��d�)|]��A����Υ�A�K��d's/��dt�&0��Z�j������T5��U�qܻ%X�aG�	)�f�3��o��&���M���8�
�xW0��j�^OI��&���pjOU�8�����!��.>Ml�X5I��B�1Je�j�.�bv�)n�8L�E�g��`@���=i]ۊ{��0B�P[�
*.baԻ_��\�Pl�m��'6a��` �r̟��0HW�5�5�H���X͢c);J?T׹xY�A%��f����E����si���u]7-�Z��5PE`gT�z��|[�kHak���>mu�7@�{��M����ˉ 
�>o0����ޱ.s�˦΁�J3��i������P�����靱s�>���Fܿ99n�O��\?���P%<��A9��~��7'ҀqdsR�ĸJ��t����h�������t���:�3�6�ؤEPM���+�a��$|<u�V(�F��#b����P��nOf�N�F^nޫMP�]x�|b2��R$>3������`T.�j�؁���9\
�;�R%d�﷨�6A�]D��fә��i�k=�,�+��AΉE�������%Y�[g�!4ľ+b����)��g��2(��8����o��'�D!�����r�&������}�L���9�����T��
�EE3��ϖ�n��@f���l��\Mh)�&W�x�B���+����-�[�F��]�A�<���0]��
���`v��"<K�..����0�>Ζ��O�1��Ê��q"������S��3L`�y�Q8dh�@[o�4��+*�v Wu�=j1�s������]�j�o�6���>3�R3]ł-����Q�fqWX�?��\8fU��R��]�(�1���g`��s��P[�H�L����Wjp�`|̌8��F.���=�3�d.bt�iS���Oyɗ8G� ��j��@V�%<-�j䇥<r�D�2PJ��TS.iY���8��&LH���E�&�a;%-o��L��a�On�-��UK�`����Ɇ�%k��R�z+Ag�"��Q�&x�+T�h��_�b:@lKk̷�Ơѡ��
�W��i;GCE@��
laC�����v�/��h�����(�(e_C�����^�q�.-���(��x�7u�����}��RQ���jѾ��,PD�~Lw��DE~�AԄ�a�`!��BCu�FB�<�/�n�$����u��Z�Kijm\��g<���
��#�Y�O@��2U�o��z{S�߃x�c��]�[�,o
����h��k� ���\7�i�2�@P��t��f�E��)D/�!�'����  �v4)�@��q�L���ѬR��p�W ��T=��̴`z���	��;v�D���2��j�!�m�&gT��9��BSW�*�9K�K�<(/V�b��D�*C��7���%;�Ǹ��a�`A�ZloMM�Ӹ��;z�S�b7��)Hs޲H!�4P�j^GT[�3Rs BeU�����:ϕp�d�͞"���OzD5>B:��,�3��/e��H3��0�F�M�W����Է�Qnc�g��8�,�O�%�����)�#���-��PgGy$k��Ex�Е�0z��ōb�\-��(�D���<O5��^�[�w	��