XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���<I�%�N�ܐŃ/��9{�oT�|eǍ#zKx��W6�\j�a�7v�- ���o�>���D��5D�gq8�)a�`=����9�~�e�Qx���"p���hغ�| `U���q�����"�ǏT'�$�a�b���g��v��V��u�i��������O?j��9%p��@��Z�	���àB�aX),��w`�{�
M-R�&�Ʀ>���6���j�5<P�p�9�.��^��Ӑ()���\@�����{����ꀻw$B|c5��G@��p�$^�/�^�'�au\,5$=��oSޛ��E����9��E9Y��i���w����Id1$�&���iʼ�����w�>���#0z�f����I��m��缍6�X��g�ڱ!����<jVs1���K�x�>l��HvT��*̲<f-�4����1B �0�T}�]�T�@��u+|e_���s�:�'g)y�1R��~B����2 ��|����;|I�����sqbգ�M(�"�����-��f����=�p;�,
����yF�!�H��Rl1hgio��ȅpF�I���J�͹�������pPK����_�_��}�p�1��J��$��C%mq�H<�8$m�|�u���1��<�
�t�A�������������-��s�	�cMi�&�dز/P�=g]%�~i������5�_�A ݴ~/"7/�v�L�/�
d	6�2�m�:ʻ.Vs	���1aM�S�)����芞䜹FT�3Q�}&ⵥӞ%լ����XlxVHYEB    b087    2540;B�SSt=i0��i��_��qfc��6ª��L�E��V�)�x������v�ڪ_ݪ��! s�"���wU������W���bW=�\P��g!rv�/�S��ꢇ�5�s�yD:T[?�ɇ�.���,k�V)�D�j�w�#��;���m��g��� �[�sg\j<'��/�������,7�\J� I�:��:AR5dK��P����ik�#lr���2$ȮD���Ȯ`y5�*�<H�.�(��-�꘸^�Wk\���M���9�~�8�!'�{�XD��Ox9���2��Z���oTpt�n�2�����C�D�R�"u ��G. f)�E�7.�zC��\=����r!n�
��"_k0������D��?3F�c�I�aK�FT�aR�1ݱw"�͸�z�Kٵ�\{��/@$LK�+��V��'��	����'� bUC���/���f7G�	8�
�����-9 ��?���`�Q��?Y�n|���v�"J�>�Ƌ����5�}Lwr"�<�s�m$4�LZ��<�Er`�RުP�Pk�6z�?KQ�$p-�Q�}i�Yt����i�1���|�ҿ�J� H`�D{Rz�qh�/�P���ɲR��U|)�^ؔ�ˀ�����z���D�q�!��<$�� �iD$V!�6l�f=��j[׭)
3_�;�-�^)��ˈ��/�~^[��F.��:i� �U�S(IiV��\d��_^Vu�xM��SN��̐R���86�U��g��z�3E�E9���Z�}xw����!��׋@քS�08:	b-�S_��/:=|!d;��c��z�AqN�p~>�7y��Š�VHt�>�b�:)ϼ<�\�;�O�ܚ�
G&��G<8n^���\%����0b�X�X��ʰ�-�#Xu*+ˑ?愴��m�](����ȠG��OO���k�c,߫�Bwͱ��}���XY����H��/#^,�/s/Y6����e�,��9C=�m2R<�aZ�~�h{���"���S�t*���%�ϛr%��|��i�?��Bg������f4�|�û�"IB�ۼ��x�{@�s+����Ξ���/�mn��zc��ۖ?1a����K��8Ϋk;Ln����G�-j���Я�7Sc��h��(f�יɪ��?qx���+� �����ޖ�V8#|��ꪏ�QG�08�݅�b�n���Ȥb�;�ْ�����F�V�r��:r2�B��(�Ň�I�]�
�G�r�F�MC�جCi���]G.�-Qu�E ��O����)p��¬!�m]*d�$��h
���a,LhI�ç�V��MԮ:t�q�[i�J܈F�D���|�t�1Z�E��>t0��8�t�/���>���(�CB�S�\�}��@�R�ASG\��S�����9a���?ر����z_���3�BT�[���j����N���lD�+�YYL��� ���wI��,})�3O<T
́pMTFUq�y=�M8���N���j�z�m��[�4��DoIP�퀰��E4)��0PM%W+$ji{Wo%r��CW�8�۠d�Wc�vg�%F���|G��QG.#���_��ݦ5���� ���z�H��Fo��d8m���hq���d듷�CR��*h��5S��SYz���s�Q#�1�\lC{$d�ة���ߩ�á�L�y��a��1�ğ�/W��L�}��߲Y.I5�if=�/�@�CKe����,�G��P��=t����(j������w�̃h���\��+(�=�^��W�_Ou��F�g�ru��RX�YQ�,Ƿ��s����<�tZ��I��U8��_7u��"FH2ya�G�\[����7�y��O+�����4���WbE]) e�Z��e�!�KR�3�u����(
�O�XpvwdA���Cu ���?}Ka5r���'k��A�d�K�����2*�q��b�L0�P�d�^Z�E��h�+�)J��	���t���$�Ty��ŭv3x���ޢ;���:6��l�%i���о�k�´c{��N�n�V�>|���f3�G�������+]T@���D%���!r|&`[��*x�=���1x? FFy/��kf�,I�A�5_���g`���^�iV�Ym	�yGw������)�q{o���jl�O�ML�|
?]��oU
��^6�����_���ǡ|�bgf0�}�~�����_W��A�6���[a��1�]�-o�׍��ܚ.b>ZC��nd�� ����!ͱ;��-N1�ϤKB��S`����q)�"���[=)<Y�ĭZ`�"#�����r���ub�}�Hb�g�ͼ$<�����l�")W�QC4&�pzpNvŐ�eؾ��t���UR
Ux����$���N� 	����bm*6g^���_���KQV�
a:�r��R���N�)O������ ��P˳Cp�h���":����Hgg��z:K\�t�WŊ�;$^0����b�� G��ih	o������m%-/�b���?�`$0z�'��q$���>.ֱn�e >
����ҫ�/!���x���ʋ��iR��8He#^%����o��?O��y̺@/-ܠ�ŅD��]{=1[��&��aɲ{�|�֙�ٞ.�H��'ҡ��G��"p��3��s�1��pT�X}��r�8���s���̩��=��N�D-xs��D|�%��P�@��NZ	��6���?��nk��Z]a�U(��1��*�+�v�5� SR�d/&�H�Ŋ�}���N!�nI�d�Vc��(cyb�*Ek��_���UBN��鰿gS��V���>�g2&��#E���\"
��_adp��"�#�Y��f�4[�z'��Kc��dф�U,<^I��HJd�4��OU�'��!y$G>�,�iM��mB��%�4Kk:�a���Zv�k^�H�F.���'�<�W'vWw����:���}�~{ m�DP�i�u���x/Ń���@� ���|�5�%����L�(�R�?�m^r�$�D@��dI�ʗ!ʆG���E�8��.�d�`����?�xƿ4��E�B�q"O��{S{p׍k\�(��%�7��IΘq�#B4\�7�-�䭡VU��Y���p3A�O��|�k#sڹs��i`�ǉZ�.l0x-c�Y�N��z6��!7"�-��dN�h*��JM��M>�h�4Ӂ��<��К:���!�*l�_�DskVg�D�/h���踀�w��<j��Ho��q�X�s�.��ŕo9�S(����A�:�T��n��t���L����ALo�\>�.m��Vк����l����a}���s(��o���2���'�e�ɫp=�5�+aO%h��Q��j��G�/y��p�0)�Q)�QfyH�g)v�DOE����#4���`*���:C�� �0�Œ��
'>��d�>-��Q@�v9�Ɠ�y�n�4��T����Ih��v�l����C��A�EM�h�[�CWF
��RI�7����94��G�IP9 %A�a0��]�Tޣ�	/#J�jJ�Ovpt��l{;>���Ҧ����u�\ 
�"�Ez�_cK�xl��I7X��ȏ�[�qO4�y���#%��hs��Dz/�䃁�Ӆ�h<ax��c�}���͊�]����������c�(�U��t����� �d�Sʿ�4��~��)�#�pL�3}�y���BIY$25�Vw�Y@�ױA�>$
���E����L���� �J�T�/L;�g#�=�OV��m�l��&�ɢN�m:��u�f�!��վ��b���gDo���L�XQ�F[@�3
�]y𧄕"�[h4k{#�$Z�? ޗ,�<�g����/1ߘ�P<�M��EȀۧ�����~�� T��?��Z�r��V�2i�j�]mŰ�$1��>�.�a��<B�'�/������-��4����z�wT+��͈�����$dڠE�~W6��G�l}D��V
�f^_@ˢ��"q]��'���<r�a�Ûu>�dP��1�e��W�}ـ��K;��܁�?v�?X�/��slQ&��_��k���&#:�r2�W��>G�:�Ӗ���d�����1�"�"4q`�=Y��k�Z�~���xdܤ�1����_.j9�6�\J'�6 �`�	q�6I���_V�/�e0b�T�d������@��V�ӑ��ܝ�/�5�#�z���Ԝ�\!�{�1��ctca��+~9��q���KS]R���,f�0<x��T��|ׇ�x�&��M��:�Q�O����M}x3¤�z��J�P���fj�%�38b �]�������L��{h�Hv���w�t\�c��/�I:��ޏh\/�Ƨ}�5��>�έ-:���>����2u���\�R����d�؄�y�"�ﴓ�55��T8�!k���?Զ��̐�Z]�y=��j
T�9����N��._�L�ԟ��U�7Iȇ�x�ye�<�Y54��c#3�-�P���@s�T������18NTͪ�h�[J(*������q׻&1 ��W�r!W����$�x��V9A;8O�D��	��y���OY�:�l���Ky9�V S�Ig��������#�(
����G���>����Ou��G�yj�r��!ϫf\�}�Ρ�n�����m�rB
̱���g���E֠A,��T�-^\���wEK��"u���0�U����:꠸��N���޵t���������lQ#��Z3�o�Ewӊů#��oq9j#[��H��o�1����q�U2�W�XQ�Q�$��;���@�NT�G~�	_�h ����i�@��\s��я3��H�N�''Uꕁ_c�pP�;�"�~��U�%�R��["7�����T�z5�<�eM`Cv����f�^e��ߨn'����7f�,�j6�ᝌ��ąJ�KE�L��;�4]V�66�&����L����y�1�!7 ����l�ڂ�Ao/��m����1�E�!é�6D'��ނ�a�X�f�
U:.��F �~X�>��B�Թ�3�͟}��.�R��o}�	���㫶:%�hŭLG/�S4�H}���Q,"T��l?�T"��9�����9���ޝJ����Q~U�%�A �6�2���9�wF�Xd��������,˯a���=�K#�H��9�⸥���JDh�چg���&�}L�;�}�>�/��*����>�����1��j��!N��N����FM<J�>I'�=V~��#O=bp��c���r���L��",
m�?�F&onre���K������O��8�a����+�Z1���f��P�!���g,����0��|F%�
��pk�đl�SEVl}z9dcL�{��T��Y��,��X8��Ǌ�2���k��O %���X�b6z�̮��S�`�M<�B?be����"͘��w~�=~uZ%hU���m��`g�9��	�U)#(��#��v�Z����N`�PFg�o��s����A�����kZ7jEiJ[�� /��B��F|�U�{��ᄧ��i�5��p�aj�r���k���o]���j�jeOl)p�jwE�f\�꿿@w����Kb�����S�����.�X�ˢ��/�L��x��F<�ʱ����LA���H�s �m��^��|�^�r�0��#����ߏ�;� ��y5k-OGؚە|��12��R�����$[1��5�9�{�#�D����
=3˄'�z�9�w�=#o�w�C�F��'����l��հ쥉@H��W�����N��?q���B�!��U�y�Z���e��5s̿?:�j��(�q\
!@���X��J�A 1�3�h�D�U�Эx���]���!q��W������B{����MZs�z	�؊�-�SOi���3�ó7y2^
 G����ӾH)^��5I�X��S�~jL,����]tsK@E����$*s]x��pM���i�o��ǟ�IS�Q�	��;9�g#E`��#[9֒L%��u���_�s�,7��???���ґ��ߢ�ʇq��=ˆ�҄ꄮQZ�Z����֣��mR�7g,�ZO��ߐk�AW�c�9�5u %��_s�qF�D��e�ݴf�*@�n1�\ �7?��9��\�$����*_�*��ѧNOe���o�͋Ȥekf�Q3k�WPa:����bh.>�kL�.lyš�X�'+��hv
�N%���ȆC�)� ȥ���"�J�hI ;��y��I��4��mF�������K��7'C|�O�r��p{F�f	��5�#��sT��$C�4\�,�2q��b���e���dn6B��%Y�Ȩ_w�+���*[�z�g�&�gS�jLE��j�?�V����^l.Ls=:�è��z������}P����5��%N��R�Z�Pf\��H���S�[� �e�f�	R�����3H�e���	^&�.��hZ|jP�[��W��l�Q�/�28���Yi��x�m�����9$-	}!�ľĕ����kE<A`כ(I��fs�U3;��&��W�y�Js�x���-ɦ8���kr|ft��L�[�����������MǵV��˖��h��QJ['��WN~щpR|����T�x���a-m�.�ӕ�9������S�rǯ�w�Υ��)��E��p!H�	��0� nz'���V��l��ӊ�ʒ��a�0o6^��1^7���~�G[ό*H�r��#�-?� ����yV���#t���N��k���G����3)8���T�a��a�#)i�#�=͝���ͽ�w�]^�2�*(�c����`h˰U6�'i�6GiWy8��d���z��5��9�.��{����r99B	��i�	���5c�Oy�@kn����ذ��5�x�-T��������=r�#$��� �r���~#3a��D���f�Z9�|����� 8�ȿ���%��m#��#>�	7�J��Y���%�qeZ���|�o~�K���D'X�@�W.f� ��u,Gm�tq�%�˲�T�wza�t�Y���)o�lO D 黓�r�TSXtQ����� �q�,v�{5O�a�PG���'쑣�tÚ����	
�)N��5`f�gy�����x<܎�����[�ۀ�X���F�34�<��@�2��?���Uw��y�J���Å�X�Ym�w�u�Nѐ���0�N�{�s�T���@ 
Cl5�Ŵ%y�ʾ=���v�gJ*6�X0-�����yq�#��4�<ܰy6t��Ax�}�x+)�Uo��D%��%��T��']6����#��n{�:�3K-y�J�*<�	CUۗ��Ɠ�������=B�H3/�$|Ԡ�ߝU��j�";������j�#�cᦨ�b�/�@��l�n��10��Ȍ��B�z.d4S��uӯv`bn�5���f��^(����YoC�+���y��>7F�KL�ˤ �!])=���(���SO���ɥv���Π�Nփ�'�E;�Ny�Veg�ޠ|��\����5'�KR�wC�~�+�\�y�\���1c�1�vB6�~����qb�(:�P7��fpn�XE*�?�MYD�B�����y|j^� ��@�e�����./���ih#�Ν�X�䑟�fd�Z���[K����:^"�d0^����]��LJB��������x�����.���m��W.���}�_����������d>���F@Uk;�h��ݪu�̃�v{�[ɂ�&���|A!	���| i��b��@c�NEir�eǶO��xHN��/�iI\POELûAr��{���[Ԭ�L�a#����=���ń|0J��}���G69o?=�y�zs(���w��~�CQ��D��p��k��G��|�k����(�1<��aVܒ�%�v�9��s��������Жr�E�di���ο����
���n�8�Rj#��@8���ϚI?�3�i�D�yYO�+ԫ��e�8a�G�y�i��� ���C�{kl��*@U�����b}�B�7B^��W��<�f@~�W��"�O�����)������>%Ns���m��]�!Q��������0K�j��B�%H5�C&�TU+���,fJ4�H_L̾�
�P�Z��tj���sa����``$^���&%؝�/�'���Ξp~M��v�n~�*2S%��o���uD,;!�2�`v�1N�Y�a�:�g��	;�-7d"*	]����)�j�R��r9�0S�ۈ��p�a|�o��K��:�6�^�]�:����x|�z���<�^ZU��s��d���M���	4UA���1�EĢ���ŀ���dt%
+�zaOd��׊TH�J"��/����9��x]��y���HK� �{�n��Uz"����S�y	�n��<�U�E�����몾k$�S�O��r4	�*�ȷ���7Bc4Ҽ�8)�f�ñ��9�t{uN��tY��F_�me�aQ���;�-u���.^>�Oo����K{9"��]�,�-f%t�{k�{�I�ܺŕo�:Z<:3 ���x��XM��S��yP@���������s0������@��P���Ҏ[0�����+y�iȗXoχ�%���F��d$�'�Ԁ���ĝ�6D8?���!�$��:i�������F _)�2&By�2�i��7M���ԩ:!\�M�Lٴn��aF��v+}-JVk�EN:�Q�M�̑��ضwo���H�UEj������v��ϧ��h%�����eMv���@]\�� 	�Y�&-�x�J�Gמ�4�O�ć���g5!B%��I��\"g��Ô��(W��R��b�p��{����@�Y�|���WF������"Rxh��Im����3���A��q�Ģ�X�6ur�$���Rb\KЇZD����K����.��Ӕ�;>3�=�G4��E._�(
��Ƕ������_�]�
�z;�i�c.�hϛ�ڻ�Y�>+��vP����dA�ID�}"�r�����ly2��\��$�7QRS��~��!_U�#�������j�T��E�Pz��=��1��9��O�����3&sRS��9X|_�z��uT�"s��`�2�7�
�ɌS4�h�>��"(�8�G�s%X�{j�
���N9��'3�j�U(���@vG���xtr_I"��� ���������ǰ y6�O3��u)��l»G͖N�����Y�D�{��e�NR|�(n��N���q&�$�c����#I)�t��Mw�u��@�ׯ#��V��1-R���H�Ф.��E(�`�E+C��C~��R���2�u�ԙ�Pj�6��l��Ż���%0y=����Lz�