XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��L�;�
T6-�$�v��u�}����u��{�"Z�WbT}l��uc�q�̆�Igf�n/�=� ߿��(�5�֌F�ꬕl��<
�V.��g���hEH<i�)4B�?[Cm7.^�[���<�m׸��&�;=�N�P����|6x�(^�䎡
aE�DMi�ц���H�{� bl��g�㽞KK�_��&u�ۄJ���/��Y�i�l.j�I��Kh�t�EM���i� /����jQ�G5d�AMPG=w�è�|iA�r R�V�&VܜЌ)�+ԏ�c�)���j���c�D0m紌s"�e�����@z3\�h���/�μ���~�_��z���H�#�x�����"ށ��#���Id����@�n>4|�E�$e,� 0z88�"���Ђ�ۢw�TEk�YN z#�j�C�m��X_���:m�2�!A�p��G�gn��P��������ci3eK�|D��Pq� ����ˠ����/"��ibP��<L����=mdt1�N�Yޮ��&�8/���S�[M����}��r9���?#�	F��54+Բ���sT���a�I��J��L���A*!&eJ������wy*̎[�-�����d�����^���j�������(k�
��;��Rv��-�5���P�@��Aq���WrY���?�n�������߄1v��(��Z`i�y����CkC�,�ĩ���V�c�qv��V�!@8���� �yr�!��Y���;�yo>��XlxVHYEB    5cad     f00ο'� u�p!8�+�ľNV��g�pYz��$�\�{֡~�X������`q�Vװ���'��GU^���>�|���^��J^'1.9�\��9$�ć@-%�đ~k�P�xG,��,�>�w^Cq1o�,X�]DJ��T�����Q��Qmc�^��j�1�2^�����Ku��G=� �|d�D����h�j�2N?�)�������^r~����Z�[�������8x�O�rs��?<ޝ�m �s'�����ӌ0=	��q��*z*.���OH|$��C��9x7�#���k��)j*���i}���}��%�p��Y���/@�!�����d��)����:��`1�7|�[I7k񨠦�˂}
�;�^2-���l���:���[·lm)k$j�	)�E�. �3��G��������o\݉�ތ|���<@5B>���I�t�c8��HR/.N�P��nGE�r��b6؞=��ĕ��<��p>\�1�x�Ld$���s�ĥ?��C�ņ�2�s���S�#��VxW(��O2�)n�iݑ�ң������%���f?�h���Z�`���D����*T(^F����u��_V�E���m��vN�IczI+�?pQ������3��4��y�����ö_��[%����J������%u�4Q~�ۨA�g��o�#�GR��P.-XWT2y62�7��XPw�+Ǹ�@�R�7�?�y#W�&"ik*v#5M����U��6�,w���Z�`J�?+�s�<��ߵ)X�!=� �a�#��$���d�c`]��E��q���μ4P�A����L��(s7.w^=;��N��b��x���0l���)@3�r��
'���N������u�\��6�##*E:�OrH=�Gݼv$�g�`�$���$4��vJ���7���ë�A��'�=�X���"��j���	\�F�bߗ�[�Tޮ��)�OR|�O�ֹ�@�˾��<C�[�/��v;ÔЦy��k��ґ��p+���{0p}*§�`�
���"�8V����#��p\%z4�4[|� ���`�fjxgg��m2�3�� �9Yw΅��M���ze��o�5�N��}2ڀ����.�%�� �hV�B�� [�R��_��\��3��i9�>o��^2�p*���1f�_6�W����*�B!جg{��RLLVw��+���W���4���X��Ou{藒�90�`�j@�4e�oO�oG���_�X�k�)&Rs�ɔߴ���<���\VZn&���8Y��0������(@}�V���� �lޗ|˟�|jrL��I?�u�����HP��%�=$�pp�v�8h	(ew�/��i�~��Aa䀋@�✎?���6��ַ+��H�;�t��ω��;�'������sOd2� o4f���x�%���@��Uv"N�n�r���)ط�)+��c��`������Cs2�0��Sx�ҫ8E}��2��7�x��>�^��~�a?�]O��p�D�"֜^��tvj;<��y��EE�!����ά�b�-rgP�Ȋ����ᄯQ=��B[`hs熆t�����/�6��?�z�"�i�T����d��c�UQ_��w���L&��BtXX��Ķ{�-�W�N.Q#8��p���W������v ��J���kCCuk����k�?��ڥ�����̶�[�bo�o~k#�����
�m�F���'x�Z���ao���h)O�IP��ܿ.=�l6'�J3��1�����f2��/�H��rB�ʳ��z�A`K�L{!6�KU��֖��I��41�y
�_(�/������r\�y_UklRk�������d�������!���G«�Pp|��GF\H�<%M�Kӻx'�V"��o;��w�$H:#.��U���-We�B�,.Ƥ��"mS�4Z�s��4���E�*����mht�I�o3�������������W��ƌw��cdL�9�#Y�v��b@J||Afp�<��W��[Lt=:�f.��
Y�ᵓ��� ��_Pv/���<��6���jhc��q��bX��đ���r�}mt�}G}��iV��ݑ�o �r�騀Y�Z��ք��,�[$�<��Dt���N�S�&z��w ��.0"r����դ ��#bu����G��bnOpg���ʐ�9�LH�u��Ķ�r!>�p��2R��ϧ!.�`��}�����^OW���(%��O�Ϥ[���*���ph5�����j2��i?�����D�X�(r1� �8J�;��N���"��:��u�*�=N]����cx�Sa��/��F�n�F�@S��Aw��(�s�=H�]��fb�W$~K2�O��XD�t&_T���7~�%�c�{"A9�|VL��(�����%\� }�w�'�� �v��K� ���ud��b&�p�0f�n���� 6'�}K�O��ꁄ }��k�T,�	��c$��`=���ů�xU"�3��
�N�6�j��i�[�1��>�B^�3-^t�1ў\am}\�Σ���ք��	]�6���<�Е�ރ��"��)�juՒV@8��] ��cd'Vg_�z�~�������_[)���yI�w�c͇�����x�ĥ�F�ZHs���̓Ü��(c�^�N
=s�.�uxߤV�w�*d�V�����^%`g+��G���w����/��N��*!,nZY��"�z���T\b����V	e�0�� �J<�_��m�V��(������ y\��|�]�n���u�c��e�!Jdm�������B��YZ:�ڝإU2����dBX4[,��󛾇ЛG���@�MQ�щ��w'��.FA�����`���|�g�T��i���}6�ft���x�l`ZS*Ǩ*d�F 䱉x�[,\-��W����]�L0�)kC�7�����z,���/2���=(v~ʠ�_*>Y,�4]e� G	F� �+[����7���W��?t�@{R����\|T�b���G�d�A� ��� ��c�Y�d+ �ɼ;����J�L7I*XZ/�MS��H~��K��f�g����4�3��{㏗@�-
]�~��R� �q�����i�R���cJ�!�:�?>;4���ah�7ս$�@�>M�́�:
E�}��DU�D��C�"KO�1��.6�߯�/��0��d2���08��ɾ8:�,i�
&�[��ﯝ��|�jXG��>o�����(�[Ƞ�����k=Z�0�	R.�|�R��]��Y?�;�
s~F��=lJ�4�J_��	�c�����[� ��SP��&;��RI�8�����&̩�����3sXs���'[>���_���j�sb��8(�������*R<����Z����M�}����=U`�8�s+Bx��^;�͒l���`�'���(����1s(i��?��X|+��mɩcn�s?αW�G���X�E�Ώ� �������W "�~9�Ekes��\E:�8�L�b��R�Id�Bc��(;���	oL������*O%��Huʗ�W�z�U2�+���>Q�AOy�I��z��Sc�h	Dm0��j4�@�Y^��I�n�����|�I���Ae=�ׅ�5犈X����,���F�Ar��*1��ʯ��/Z��]�� C�?�-A՟�|)�*�&)����jє3	x1g~�C�h�C�ƃ,�J:�XV�D��ԗ��K�Er?�W�6I�+�"i<��l��$վJ���G�aw+6¡�+�D3�{�����&zJ