XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����gsγ�a�ٓl!��T��0��d&�_
/�۫�$��Ȓ:���a�>�����J��'�̫`j��}����Pa�a���(FQ�"�t����
�;CK,���l���H�i�΍Rt�4N�l 54q���5x7f�,�i��?�W�˻rw���������^�P��Z��W-�۝�����E�9Mh֙uf�'��e����ß�4�o�$u���+̀u�D%�h2���N:�'?k��W��Ŵ�����/���-�z����o���X�ed��S����A���1�V�C�L]Eݥf%5��r]�T3�H�X��]���pV\2�a�.iA�A��<��|��#=Q��I�Hlo�ˀLT��<���>ɡ
F6j\>�0A��˫J& h��y{\��Q�����W�xB砣"�r�I���o��6Pko�U�c׈��P����ΞLX�0�M��+�b�S�U�b� ���3�:;�F�>��;��z|��J����q�_1Q �̇�Ť+�),{*��'�b>r+(�P>����>�>��`ha�-:fo�����q�SFQ�3��Z��H��ơ���*9����>y: d����j��;��eg +����#fߧ�rt�2)�� �d�c~:��T��\g0rHr��l[��3�X�[����o��yLʿ�'s
���װ �4&�|��ؼ��mO�d�w�>wh���sKx���5#��g2��(A'�^x�]9���کXlxVHYEB    4284    1110;"m��G�������m��_̡Y�(L�@q������d�1��VdE_۵�a���P�Dpa��9�jR>�h�&��S��0��5M�����Θ��|��K�J[�]A'|��g���"� P ���O=���0�J�DV��޿����/��!�%=���K,�~�9}��Y�{5�l/Q�l���d�SHT���ʿ��v�°�#��O�^
�P'�����n�rN�����}EK�
1_�����)�Z��;�qjf�~�Å��0B����8��3õ�z(�O2�A��\ցƜ�����?'&E޸�Q͘"D�J� .� {��u�]�N���F`�`!���cO�j(z�����Z �49C!N���]�
��98�}vyYsWdi��+�G]���G��h�}E�b�^[>|�E���� 5�dS
����Zg���p�S�]=�"�Wq�{yv|F�M���ѵ�u�ntk�m�]y:��ɥ,.h^ٹmÈ��HN}I�H0C��ZG���
g0�Cmd�%?�H�X���P_�}\�2�.��(�ؘ�W�/��s��Tk �0<�?Ru��GZ���y�IA�kɽIs��6y�x���KR�l:��)V�L���8���,�q�zl��.����e�==��,	�k[�,�˧�C���t�,�Xoi,�va�cpMW8�!;�CcP�?�]�/E�8�!�0V]G�b�v�vW:������9�B�� �������c
�[�u�د��,B��,�\`p>\��޾�J y$7�)^P��d��?$��`	(顧�:�E�&�F�?ԺB��A�a�sn��+q8�b�#�s� �]��1O��z�*�� c�V�\�Ǫ5�ƪ�bw՟��c`�g���e N&����1�#vu]�O��pA#��,уK�d��2_���IZ���n�����;����:=���F�-��g Z�7��J�s�f�	B�� `�O|gl9�4�-�%1�BRú�>CЂ�o��%�aik���M-z(�H %Fc"����H�2|v�X��[��QfOMc� ğ����6>x��lZ"���B��IG�|=��֎�Fr!qYH�T�۟,�A����ҍl��U�����Q 	%r��j�:�r�}��}������wv�[[`��6ft��Ǐ��Y��@M��$�H�7�z�=o���09G�	h���$��0�d�	}HS`��5Zǽ�����
�g��5EW��qZ�](Iu�(�`�Ĩ[0�����)�m��<����!;f��ʷ�Y�TU>9�Z�z 	=!;����6ظ�OF��6�0������=x�q�B8�mhu��efX�'���s{
�❶�$m@�N�ɾ�:l�UɰKnB�u�,@�E�O�#�[J��3e���޼��	�t�<�'�k�V�"���"�륂��cBy������<{�OӅVu,�׭�� D�@Kn�.���:����LQ%�h�*K(Μ@޸�㪤����x}*x)|������C�/�M��#� RxH-	��`PEĊ��F3�yx���h�eaqm� ��f$��b�>�>иƌ5x��>�mkZ)X��L�-0����t���-uT؄��V&㊠��t��^U�ˡ�< �rRǺ��s��h9��;!����r^A4�m$�a�/p2�j�p?E�U򶪤E��r�G�)�V��p?}�]�@��  �?aZ��}{H�o6͇ˑ�?y�P#��T8��[l�Q���݋h�y�V��h $Tk%��DR 1�67�+�F�,}g�8x��X���Tf�Gk$�E3���oہpgjT�	'�V�7�pړ��I1���H}Ä��] x.���!��q������$��b����T�;��}��@�Z�0��N [�j/\' =�����D�3�[Q� ��H�D�������&�}��|�oB�S�r@>�3kY��ZN^l��hHJ�Y���EՀ[�'UAa�<��Lѓ�S��g,+A�R���9��^�~�4M�ieuf̎n�d	-�!/�v�ʲ� ���e0�T��p�bx����#�e4n���|�@d+DX�2i��L�)�7�L�u��w�����!6K�둰m!�Q����v�ѵ%5s��G���c]I͑�V���'"솞�9yUg�x�h�"��!\[�}���c��N���J��3�>J0H{s��M��4�^ �q�s�A�!��X��O Zln~L�-D#'��'� �v8B�+u֕��7��C*��`U>�QQ�u0T(ßV��|~-������|�������>��E��`K���M�����ԃ����{'�.��7<\�s]�Ş݁�kV7g$��sf�5 ��#	��_M�.��u�C�=��҂�U�j�'��m���r(�C�~�)��%�ײ�p)�Sh6J*;N@s����p���բ�'�L�.J���\į���g��ܭ�v_֎sSd�D+�aǿp��4�c�<�Ԩ�["�E)�]�BZ���D�M�NG�m��Tc����P�MT�kgҶ��pH(�Sgatއ��L*����N[����L�Y[���:����uo�))i���e��I�YON��< �ϿM��O?�p$��F�
Qf�h��ø�L������4\ｼQ �����A*���Mv�\���F��@�,TN���α��u��[w����Ήz���=v_gw'	S��<ȫif��)]���y��W<'��Z�@䥉����D(ۈpΩJ����?n�e.�T�h�;AKL�g�*"�q��csE�%��=�_-�? ���4)�ӡ�6M���bۣ6N��\��o/�z�b�j?�;G�45Y��~�������S�$�Q+Ŗay�hWTzT���q����Ǎ}wm�����Z��g���٥-z�8��ΰENO�x�F�ѷܺ%�5kCo]lv蓼%`V��l��=٨x�3��@p0X����6~��ٵN?q�눡��%A�F��%P���.�Z6�1#�2f�x:�Ex`�����ֶ��e��+�+H�K�DU)z5)�qb[϶?w�/y}?�Ǥ�HY鶞 �+Ű@��͟����u8��J�L�cn��.̓[	��Ǌ9h����	�Lw���IE�1���|:PZ�/���R��Nu�r��8�m+.��JH�Ԉ�5cTK�q:�W�_ݢ�w��S��P�Uo5c ��K���l��j�_d���v�8�R�|*:��=�X�Q�G����|��N]��q���`���]��~`�^���K�A�r��v%��?z-TU��}�������G,)ȕ��$4�����P���+䆻Eua�"��0�)n�+� �Wlwܛ�yN�.q�fg�֑�[���Hp�X�_�*}h�-X&:���w=_��1��w��v8�U�?XH�K��:��+�Jf��v�<�����v��^M�E�PPQ�?D�k�"M.'�+����Y��B��o�h�����w���}�H)5�_����p3�ơ�%M���D�z��2�^�7��K�9դ1��0,��a�׋In�����◪K6��)�L}�x3#����
��S�O�i]���@1ZRz#7����1 �h8��:f��T#�.[�����o"���[�1y�F��P~�h���f>/gv臈c���Ѐ5DHy�矈�?�N��}ڗ<��m����ȅ��]���;���.�+��b��ي?�ݞ��:��M�z���C�@����p>�5�|�D�˾����?�=֒=�@���(�l��1�֐��8\r|�"��J>�U\����{'[�����4x������X���3����߅y����Y�����5z�~�� ���5a��E�Y[�I��w����FB6�|a�gjJ�E�M'��+��C�yB��Z G�z��\MV��H�����a�*:3�r�D"��8F�&ζ��qHL`�PJ	j�x	+��pH1�)����m�i��u��j@$i��CA�+��'�1����vVC�- i]����ԑ�DL�������"�Ձ�o����"8��1z�r{��*,I�],��#8s �<ŋ
�U2P���V�J�_` ���؟+��,pV��ޛS��9�B�+u�?df�=�A�Q����G�|αM�j��%<A��(�j�4�-��2u�(2A<���	8���kᛘ��!�V�l�r�	�u>�r�1Xa����b�OС����ǷPr���G$��6��4<řE�ȥϿI�P�^n��ֈ{�d���n�G#ѕ�n2� �_�9N���矄�g+���#�ߟ