XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��^�����^��ฮ�7u���l ��w~20%2�d53�c<������`�wȰ�����������@��L�?��|ߧ:%�|p���LU�Bd~4�^�!� �J+3�=��3
+MY�X��U��]���r�ìAV�C4�O�ܯ
J
��x�HW���]���1}���O4O
�4�N"�(7��b��l�:.vgu���{ēB�_��kY�X�Ă�<�����E��>�+]�����aZg���7��g��-,�f�<R�|E�R&�c��>D�ܒ!��s5O��ߡ����{�=�	(r�ث0���M�eZj�;�S�i3I%��/T}�M�q(��A4��V�˨����*$}M��k+?9Yu8���|�v�/P�H;��.BmTa}�z�H���	\lJ���]Q}Tu@m�ڃ3A��Q�up�ӐU�5���gi"ZM�N:9T�,Sg*Fz�<��#s��ǃ)��?*gH^���D-iY�8��:�2��!�^�U���j����&^;e-�)�]\A�<E��yO1(������\T`���\V���~�����>�"���Y�KC�Vd3��T�L�*2�N�����3W�E�i��P�q�Jɐ�|
�q)�7b�UJ��V��Ѕ���ѮQ.m�9��_���]�xRa�&cC��V	+��8Fv��/��G���8�Fe��4�.�\<֘���Ǻ�B��W$0�l2]��[K�1�0���[�w�\��������1*htUHXlxVHYEB    3e93    10b0�ا�l�8,�u�ʩpC+ T�kҾ�7��$d��J�R��o�"A9����ž,�:�1eR�
�J�^ԩNm	L�����6d�����w�9�M���L�J��FrSyğ��9�Ʋ}�?�|�I�+9�0���%�� p�_��z�bo")�>���23�|�!��=���z&^���[�h`޷���(RJr��]A۲*���Y���H[u��P����e�/A�Ԣ:4�`U�m,� ���7�Y�L���R�J�-�߉�t������Y�T�O3�:I�e����7Q��F�B�ʣ�+}� ��w����� �m]�F~�^���OS����Y�����q�E!L�hqdG�V}�0S4]rݯ��<I�R"�CG�� ��g��ێ G_��c�rE��q9	5,��}��>©���Z�G��ME>�!�w��軠����)Q�oV^"���k��,�?�_��u<0�|A��:�l;�Q�J���Ӻl���r*)�.�Y>��_==?�y�j���v���H<蓖�"P��}ھy���� ݲ�-3N��:�Db;�{���;��!��.�=e���O���ʾ���I���ʖ�rRAe?\����WU��w���-g�g��J��\�k��v[�Q{Rsʺ/|��ȳ�V�q���{��������o�$����D�I�/i&\��/�Qh�!\�_I��3\�A0gu��gK��|_/�[�_���<�z�f�OSb���T1([�p�����>��^��~60U��
Ț#o�
e‪z5��1#l�x������Ǡ1�z�tz��ˎ���E�-�����,Hq����=/�-Xh��g�ˇ�n\#m/�?<��a2]}�mx��|�(�ݔ�](�<,d��:����I���n!3h����j�8���(���O
9p[�Nn�.����PHpi�����M �Q�G>zLF��{b/�pQ���QK6�K�8>J6S=j�' ŗ}�H�Ҫ��ѣ���T��2�=�ZB�����(�O�x9,
-�!Ih�w�F"�Ŧ�$�_�~����u�	�25�jY�u&ӗl
����������	�ǟx���t��k��F�Be5У90�v᷻��c�I��*P���e��c��g'O��B��x?.�ҕ���Б}t'SV�N�%Q�3��uh^H%���:lF����l <m���X��{�zw1p�y��ܐ��%�K��igUwc�Xh�V�P�>'�V%ʒ��~Q����c����X�Tj�HE�\U�w;�
:�c��܃��knC�N�m�g���J��#םh��zX�dY2A5Gf4X'��P\�c��NX&4p���7�VQ�0s�P�9k����$��t���3;��J!Gq[w�ů7��.�$�iTW�mFQ�<��I��Tb�x1�s�7��X|�U��$}T�����J�>T\��D����v)9$(�UP!�G����j�w���U�
\m����4��GE�����B^�פ˒�t�7;�O�������\Y�Be��/ ���b�?�a��(� ���ҽ��v�(KG���m�m!ݏ۠z) ��#���������N�OkS�mD���펧E�Lɭ:l0�ԧ�N�8��n��[m�6I�*�>XڙyX�����80����3��:���?˙&>�bD_K�ͺP��E���Hb�"E@��x;����ΫJ�{�[t4
�á��~$��>KJ�����Q���{��JJ��1��	�%���u�2�*J��]���s�
E �v.��Z�$r}��c���2wj#�A뭾d����vN�qg{,�/sMۗ�RτA� {i +����:�gs�tIi�������,���P���뤆��&M���dR��������ȿ�fk̒���_���އ'��獪���ᔒ�Qe�O�s�������XHq�S�T���B;�Ml
��( ?O�����a�$�,;|�d�7}
�������kbt�1�.�C�?Q*�X���k�RФ.JA��]
Sǯ���-\�>=�k����R<���
��[�G'��v �=������QE��:%  ��~{��^��G{�@�a�EK��4g9��{�@O��o���,32�g=Ӿ܏t��:�5�*��כ�ݣX�*��^��jm�h���2����/	ӓ ���D�Ԯx�}�$_��K�:��Ѻ�<��,�?.��1�	iʤj�;ĝ&�BŤ+�#��h��<��uYx�P�^����=�&;� o����.���A���+a{�4�0�֣m�+�*n�D��%����&��E�Ⳣ�P�R�eJ��`��Lw���ʓz��I���w�iɢa4SEy[=?��{�H�lrC��*.]�i�oH�Y5 Y��vЏ�/�0���N!盵�s�4�9a��CQd
Di�x�	ϋ/Bo�\FS�l�v��y$� ����˱�:1ɫ;�/�#G���"U��űۑo�pK������J��Vb�t��lM���0�;��-�?|�U�[���0���@��1�p��r�,�eV�&�5����y;�(�fe��e�ͼ=���˙�
(PS��E����ӑ�I3�i��ؿ �~���^Hc�lt�]�ǟ��S���k�8����w�-���1x��ˢ�1�f�`I�0�`{�i���D��?h���V�a�$A��S�W�T�-JNHG�{��8om�"�^�S4[�ZC�nE�v���>1(���Y7���]����DrN���ӚW�j(���>0s�!��P���2H[�?R,�u��o%͎�tb�$qNJ��F��c����wM�=9�}�c�� ��\dL��ƕ����n�)�]��~�����P!3�混6�?r"a+:NQP�9��ya�MBz?�N�h�`�:�ɟ�WWB<�/xt�2D=�Q�H'��}ڎ��͆��S�
�I2K�Ѣ��1�r{��m;2��ר����ST����^�����_���B���4��e$��0E3$=5w/Mx�[P�k}�]��r�3"��S�PDwhؠ�7�T��]C�lLi5���I���dYֽ��q2�R*%!A����1߈������ ���y`ގj:&x���M�]�L��\�B�����kԝ�~yvN����#������v�7���j2e�q�Ռ ����`O��t�Hj�Q,	l�2�IG=3}����(�P'_�<�A�M��i��$���a!�h3��᪃�R��`�{���Ĝ�2��%z�Ve�>�OxcNP7g�zĆ���M�t���Rݪ_.0��,�����b���{*��h]�.K��R�IS���K��ņ��$3pu��zP��9��r0���33�|g�I����klW�r��qK�#LK7�O�'���P�%3|ڲ='�
pA�1�+^š%Pl���8Pk��p��|H<Ѕ��u�ۜ�-JHH~��$O�oP:
��>�|΄������������=�_�!�R�ɾ�!6n���Y�1���1> �SvF����l�,T���p��	O�m��S���Kw�A�vq@oL��(J�y\Q��Q�j��C�Ri �X����a����q�(�!<�5^:;R��_Y�E�C�N-J��$u����4V�q�.O!��A���q'���7y&.dkw�����S�I����2�r��S�Y�۵g��ڢц��	n�)jR�v%��KXf�{sg���/�i�?����A���..l�rk����:ϒ�ޛm�����=�{�b����ɂg��-p;�$�?��l{�c̿Q���2�/p���}ݯ�O9�vְ��?�I�!�@k��͘WJb�*�_Iٟ�4Na���[��Q6��k���̥��/���C�z$
ס�?�p�n5�����d�ܳ���:@�i`Q�ȓY����wf�Aa��VAB�H �a�"���\рRYjbf}R&4�������D�^�"��F��,��;��`6'���w]ڋ�M�[30�@`��E�k�Y��@��i� R�'!Z���0hܩ�,%G}<��Pװ���{��i9U�y���uQTe9jZ�$���}��Q��L�-�@�S�f���v.B����\ju�>��I�Z{�d'0�u߅;HAYй�}�$�_�g��Vc{��Z���\�����u�y���}��5y2��PVRaG�l�