XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����I�)��$@��$���{L�J%�B�'�7���~�2�� �.�;m��A�:�Ժ�?��.�q��� w���,���'�E���.�P�/y��- �|��Zq�*��o�>� 
'��]8k2ɼ���3L�7��d�u�f��������FĹ�a%x0q*�����lj��~A褲A��`�4�ӌ����_�S�d� ����_+�t��'YŒ" ��Ɉ[9��qh����w�o�����&<���Aچ�<P��zk�鶎!�U.i�Z��H��R�����n��p�*��85�}Aڞe���|�����@}q?�l���cB��Ba���z���n��~���c{�\X#�b��'�U�|�4�9D�/��n��tJ5}��^��5<�D�:������m�t��1v�moE����9�PLY�����̉Ł�d��O���0� pg2��6�q
j�ܱ�̗�uƝ�ŷ�^�J�s�T�K�U>�y���@����wCs��#�K�|ە�%�~��0�u`��M���c��́�����4��?u�0!C w���5.�v�u��G�Z�Izx��]\��I�>U�8W ��a��C�]�+.�*�Ԍb���J�F��3Rri�5�������&���"��QiA9�^B&Ԥa%5��i���ή�Fܹ���9�fw�Y�Ly�H�ه�=WZ	t��H�өυ�ȣ·���|�W����M'�Rw�0*F��R:�UQa����a���.p P"v,U5 �}6���J��K�Y��щ^XlxVHYEB    48e3     e00Mz;L���&� +��2A�'�by��ZT��i<���tfuQ��x4u�F:y>BO����̅��}Ԓ�FT�QS�[U��ex�w�!�9G��n�?c{�;��,�E�8�!W%�+�I.�A�Ĩ���8�����h~uW���ˮ� ^���ӫH�	�kSy��Lz�_i��,$�q�$}k��l���n�V�\&	S�ϣ��_��]c�]p�$o��������7�=�*l4����Z��Oq�z�#��K-�����>��9�\W5���ڎM�"�h�=u1,CV��غ���z�S���I�8\XJ����-�p+ѣ�g�Z�N[ZLe+W��X����GՃo5���/6�Z���3:%�E���V�V@rC�R�D�
�<�#��à�Y�迢��;�Q*?�MS3�(LC~8h������ε��L������K(?C��9���7Ą�/��<��<��(�[]u�Fs�́��Tl��ٗ�ְTsЏ����A�$�{k:V�����j�&��D�[D�1�����Ȳy�.�<�pU��u�/�4�Jf�x3(;��U��b]��d"�|��I+D�L�{F�$�NuHs��Uы
߲�̧�b��Ś~$��h*m�;�����rQ�ٌ+�}�s��f܆����3pT9!��4I�+����$��2�&Bq����z���ᆸ�x��H�����&�n�BNA�Mb�m��R4��T=PzW�ʲl8��c�~b�߀ßg+��¦ښ7Ǯ0���}?�e �������u������ .�M��x��^K�Pچa���܄��eP��aiް�wM:�2g�%�����p���p4z3��'��RY����*�	"��t�;��5�X����DxvZŶI��C�,���Ȗ&���y��ʇ4��Ѫ��{��}l!�{y�v��Tצ��xB�H��"��'Ǿd���TJI���ӢY<`?3ܑ����Y�n��{�l�7ȱ��<�E��As,��� i!a��R��
���n��5��R6W�cT�l�I�lqMy#%��͞�#�7���9#�ͱ�j��vVp�H�
Ċ�3^���Q���r�	iP�[�up�W�
�M�QQ^�L=U�?LX;%/X��]ˊ�+��l�J��3�Ib�,٭\�;�D~3?������򔘙
o�� ՝��m�����׻V�Qvm���;5�z�zV������4(����J������i��ˊq������:}s8��"cr�9��G��_��>G���J�zmoaP��hd�ٗ�;
c�nx�=��q{V���ؼ�F�ig�LbV80b�d�yv,VC�YX5}����i���sB�~<�F(�6	���|O�n�O��
Ko���q�>q�"z!�KF���,�pZ����l>2Z��-8,e�b����ǲ5@Sj�-����k���D���w6�dF��R�
��'�G�^1'�.66���S	#W?O��i�i�7\����x��j�/��ֶ��q��K�qt���l�%�u*�M=;?��<	��DB&�����5�Ϝ�2��t�b�dM�!8\�R3"���ʼ���zz��]�fZDA?��ʦ�w�ůwp�qn�?��w�Įu	�H�Yzt2X��E ��=?ğ�U�o������Y] l0������T����9P��;��JlC�5�����r�a�{e?�;D:R}���o{�7VA��dXG31�*(4�;���;�M
'�]����WqjgZ��W�9�n�~f"v��$�"�m��N���{���d�	�I����L��k(�s��g8?�e+�ü��t��^�2ҍ��w*�f��K�Qc�ң�[�A�Xc�9.�B?V��OQ��R6��^���H<a�#=�+&����1Ws���е��Mȸ��)�߆���;	W��|t:�C`��K��ח�0e	���G8�%d찦,cݾ��V�F�-�zۥ1\!n�>�k��� ������������5	�1E�e��w��ɽ'����q�?�58������Q���^2٢]lvoY��)�^����'_���h��z���D1|~�y���d���d\5���b����;���V�!�1�_V�1j�*��L��t^���D��DvȤ�t2�5399��Hwp�tCo��Q�&?ʹ�])��^� #�嗍�EޕLJ� E:�3k��2+)��ֆB9l�w�L�Td�F�濖�<�ꭶ!��
�	�M�OS@�ɝp�Ol�������ߠ4tBG��
>$i�1�
��Fgb?=��NKD�I��=9�ԛH��6`���7(S��h������^�}C��M���A��M�fW�ռy��gs�t��`�M�76/���m?Y�#�1�H�?���9KRp��O}J-�S�J�`�/�mB�+z˧ h|<:�?�jېQ��N�Y��jM?��xv�!@2/-���_�R�B	uDqqw)Б��
��`&ż�Ũ��_���Qf�H�"��1u��20�α��luD�M�j�t��C�ܮ>�YoW�7q��W��ռ�|8x%�AzV9}�t�d��Q^,���� r��F��c���������K�X�[�v�����B���!NS�yM�X�,��9t�g"W6���j2M�8wt��'-�g,ܽ�܍�,*>rsǾ1ۈ����e�K2k����k�:6�j�k2���o�̠�F�i��J��і u���1%}�~2у=�2�p�L/m��@����qF�%�#`��S�ʋ$����ER]͉8�f;�b�l>�(�2���1�_��u�=J���Aq���#Ʌ{L�ʗrƈ7�g-��4�C�V={��Kz8:�_�k��6�~�(�r�5M�A31�?t(JG���HjD�Q�Ӷ!lA��5p�R*��Q��F��U@�CEu�E�#��<��g���@u�I�ߍ�eX'�M�J���`x�@����O���W��R*�1��i1#����?8��+�P�bٕ�h0�!� Z�gQ{��,�rx$�lwټ���W�v(���j����l��l�g9삲�Ra���������2��)�#���ϑG��E
=ئ�ZZ�o�<�M_����(�|a#�]��e=m�_Dbd�)���_�!\�?����ב��7',˄�f;�Uw{�#�8CY9����5n�{�h����@��4I�`T��ƇЁTϷ[Z�{(��;
���A�?P�ʜaxT&�8�v��%�I��e.��@�T�I���Q����9�2��+�I��9��0�����>����%��:LeԕX��;���fqT��T��1������E�N�E'*�xG����M����։���'�=�!p+��n��&����#�~����
��b�Į�ݤ�4�;�tA�k�|,�H�;��OV}|zr����Y�:�l{KO[����!����M��������w�:�=fO�F����[�9Uw(�����
{�N���/�6f��T!��8�k=7��:{�A����4a��#~EF�.y�{G./PdTH��Z_�'��+K/�M5wUA�wk1��[�cvk�&�݆%�