XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��2�W[or�?dT�+��W-Wt{Wz���'�����	!2�z�c��/,�W��0�8.t�b
DT�/�x���}����� ���"��l��ݾ�f�gAN�#�3�Z�aE�@�|��u�skk��? ���zC�+�w}�a���^��q\��A�� ]&��&'	~1b�T;Ş0'#�<�x���*a�r�{g$���00��5J��|��{6�$���OvU�
a��S������f���
bb�|�!����_�6�`�n4���:)�N=��9�Y�ov�5
^9
@�b:ɍ�tQ,gg�����1?kD�W�c�}�9;+q�2 ��X�;	�]������ <�)�� ��ݯY�į@T!�S5�pFS�]��#�.*�����VF�BRy/���՟��0E����%=�S�o�oR����8�m�:q�"�l0�4��Q|�բ�ESF{���'%2-�� �v�Ȥ�T�z�v�1��).�6����#�$ZX�,�m����G��°��� ���[㰕�ӕ��c$%��2��o��m�&�*�*� W������r�'����1�؜@��O
�pP���h/�7sW��gYp�2�ͺw�-����o��V�C�?�w�.�mu��.�<d3Aѯ�rFD��2ϛa�' ��d�:mrQt�f׹?��'�Z������{N7o��J�Ɨ�-�;�c9d�:���gR��p1ɤPYW��c/��-ƍ�:�q��0����*�dh�.Xs�=�Sl�1�XlxVHYEB    2b39     b10����$���p�d��W���W�i�'���%���]����x, U�L�L)1�;�?ߪ�����D>5G��
�4HKG���6y�� ���nRhT��W̦[2�xB6Tە��'�@)̆Έ׿�׭�XZ������?�,Z����_��E�^Y �HN�D�����!�x�u��H|�4�F��Eŏϓ�$�z��=%�[��߻�����YJlӀ}V�����t��}MOq)#q��>xA�I��3�"����kz]ڶrv�`�s�ET�Z�u��j֥d?��7�&�hY��<�_��\85Į4w�g�A����nX	��##%��:��Bm�#8��������[�[?��ߛ�@�w?�|r9�
�6���O�<��Jͣʰg�bx���qb?B,]���`r}���6P�j�@���������9�?��7�du?ŅN�ޙK��4�|���f('|=[�%��At�{^�Βt`a$Ac���p��?��H�	M�~��h���!ਏ�W�Ϯ0kG4�B~��
��Q�'6)⠣9�͌b�޿��zZx")����(�H��b5��ُ�h׈~v��\����j���X�����I�u�S�����^�SO�vlN���G��<'q�̘�~�E�I)
�$U�g�ؑ�&�o?�:wIFy"k�v���D��ݤ5v�����V��-�.�BU��6�O(r��ԛ뢠:W�ƈI�EUϔ��?.�Tr��G��)�'&��8w�� ś4e�3�\�
6@[e�l�'<�!.no�7h"��h��v��:]�t��6�����<B�4eg��s����?#����:@a�^�1H�ֵt,�xjs�y;e8�lo�o��A5H�vT|WH/zNz��. �R�ep�S��&MZ� D�qEζl�5�pr+���B1����q5��:u�%��D�?z��B��<#qd����_Ym#v)��l�ںB13��O�b���g�EPo����%�M�s��K4^���Q;%��t]1�����:���d��Q��.'2�H���C;�QDR<��}�NX�D(/M,��W`��'�G� �_:H%0Z���I��m��P�	`h�ޟ�S"�" 6��q��Rn�AT��5{p��d���񸎻^,.�Gq�r��7œN�������U�\�C���H�Xj�4\������������U�s��ɽ�Hň��#*�݆���a�z�:�9j��L"��5��e���#�a�bmf��{����Try�%��f�~.�X�5�UW��뗓f߄�1ԆGޚ�{ڔ꺩���Kx�9����'p��G�J���l����G�J�wؤ�`1~�mcEW��Ze|���Uꫨ���p�<A};�V;D���*2�[��z���y��	��`��j=�p�!�����K��Y|HœPr��Nr<����&=s��)�EtW�4�.��72�\�\�Z��'B56�%wX� �B�bM滢�]�>�`g9fM��(��#��Т�ݵ����om�D���#���D%Y�o����UDUClp"FV:�{�H��4��jNx�g�����+eb��OM����C�^[*�G�C��QH��G�A9��
��~��Q�뒠����"��&����Im��J.�k��CS".�| ��b���,p�[_Mf.4�D�ܭ���d$a�v��A:�qv#�7jc�&���,��������S��:���e��F�����2N�t��L{���1���c����!�,���1�n�Βs����n(LV����K�
J��`G^B8UT·Ex����T��ZF�N���SJj�����%e�>�R.p2�v�;	�q��I)o�M�3c��\)y��^Q���|��͐�Ӂ��W��_�P�,���"� ����q	��M�ۥ(�vз��'��Zq]�X*�[04��U�[�츍U2 'GYvʖ��۝5UA�L��؆Q:?_mK3�n ��u�mWju������q�ON�f,�D�㻳�s�ki����������H"N�5Lۗ����5��l1ԠKH�3�x�\;___;���C�.�+�R�����e^ݣ\�r3�X�J׸��g��b���p��͹��@S�48?��JӼR����e���o2���"wh����K��~�3O��?	�5�rw=ey��w(7��}"�߶���c�)d�-�Q���w����+R���"<U��3|�=0f�gv	^f�� �'0��°5�T3?�3 �'��<�]������̷�j����FX@�
t�EV4 ��B��\e���gŷ�(��|4fX�Q�;��P���NB���Z�����1�dP'�F9�7�-�Q�����p<�g�X�_D���.9��qM�Co-3c���c^THbl�̵���.���P���o�C�/���$�2_G=�C��9&�Pa�������R)ߛ�+�r{����{n��HLШ��B��nr�0uF2@E��}��}>��w;�i��ƌ̊�4�5}� r�NY���pd[v�0��j��p��-�����h�SA�2Z$a2
y������J4�X� �HSO��Q��1���c��Y��F�=��{h�[�k�S���a��7��'P�)'��d�E�I����~��\vhtRy�yT�
�����4�Y��D�����[?�B��jt�����a�$i��))9��Z[^;Q�����K�Aݦ���=�__%e!��,G䪢$7��P�w���Ų�#V�ωem��� ��ǜ�Q����