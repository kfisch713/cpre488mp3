XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��~�wL2X�Ɖ*9O�X���ϒ;J+K�͇¤��^��H��\}�r�$z1��$@�����޸V��Yt����6_f��D�RJ���]���߷b�}�S�~BG� +֣�1��֋�7;�� �)�,���l�NPKq��D�8�7�� j;����f��zN�u�3��@����~,z����O�����/���J���b3	���Rg�f[�]�q�Vm�yS��C�//$E��5-��w�0i��Rcg�;��^�v)0gT��{�mj��y���܇�s�fT/-Y�^r�v�S����u��2�@rO���7��A�~�_��݊���22� o�-�.[� ���L����S������W5��W�u��,V3 óz,�޾g�[i���䥾�P�����,^�8y�c��oU=mEH)��1�=qΑ�JH2�د#�Wם��v�e�����N!�x�B�Py��W+��O�:�}��J�b�;1�J��cS�ɏ >0�U�����F��~˧DL�CZ����[�z�Weg.����=�_[�qO����l�υ�}�˓�F(��Jr�fhDP	ɭx��;��"n<ќ��s�\2Za����)���o����d���2=nX��A�����ǀ��hO3�[�WW8c��v��M���T.8���rř�"͗��\.�b�ߊf��E3��F�{��{xZ/����*ϛ��vD��$Աt�0���Ygi�<������;�� �D���1XlxVHYEB    95d3    18d0� `�E+�U
l��r�mqJ�c��mJs��t�7F᥂�W��Xլ8)hE����^o��:<�:Պ��N`����E6��!��|����~D^��yz�~����G:cˌ�x6�+O�˒w�7{v�.j����}bﱔh�kA�*E=�}մ2��; � �����E]�2�����Iv�=��]�\x�;�/�����m�����'��и�Y�D7�][~Y��#�����@m�K��C���hzL�w���8��7�Sp��)���.�\x���fa��f�3-����;�4�1��0o�(kB!�d���ܓz�L�3����>�P&]-��R����u�>����o��n@�K�	��>gl�.��5�<����gsmT��g�Ly�ݙ��`0 ��/���s�^d���
I<ߤD�e���.-���\W��|��%-?x����8�ݝQS�痩������!��<Kg�b�I�s��K��ыÑ��� ���9�
��'Xii2���*�wU����Ym%�3��.�^���p��F�n�F�|5��J�9z���N�~q�e���^7+d���^!v��ߘQ�sW*����;�6$��?(l Þ��	�4behBo�8�� ~f�Z7ӵzG���	������������`�]���j;W��Q`(����p`?p�8s����w�^$y� �(�����-B\+��Q�98Pr��0v�G�o������:_��׹8>O��F�)�qXK�����k^�&�1E�A�Ub�G�w�Z�����=�r�X�yP1���)�(�z���z'�D�:|��X�.�f�;�ң��Y��G��f�F�:����g~��yr��2�P�(v�aj,ЩH;��斤K���Y2��v�����N�A�χ��Hq�Y�Ÿ䐙��i3 �����U���WC��n����� z��N&�-�7�h�h
���/�����z�~o{��B�/%����P|_g4��X>?�E`2ۘ%)�(���~���U\�.�s Kf�>y�
~3���ɤ�VwgX�h��o��	04P:��(��&�1�J~�C]#�_�b���B�;�AF�T�\\�C���	0>gt�������������`5{�}�q"�l�=1��� ���\8}гz�<)��N�^�^�\i+\"ƒ�5���4�o7s�2ɊVzSA�E,&k��L���xI?*�j[�s���Y�9S�'e�NH�͉j�I�r�m��nt�ٜU۞|RL�-x/�}w�����q��5�:n�o�C,�]o�8�k�`]�RP�_7�[�|Ԃl���a���b��\@��`F�[J�鋾򋩌�"��c�VMS�͈q`�z��;���D&_:��S�t�Օt�.K<,H�G9>�;r:�5Ȃ	-$��]�CnFf]d����^/ w�*����������6h�U�S}?�B�7�_��-�@���"���D�'��H.�<��]�_�)S4���C3��_�5��h仱�`�
T:s�
YT�Z��GW�w�����GQ;�T�[�����jYJAzЪ�U�^���eA(�cG��Wՠ
c>�0������ �t��:���.~*k�h�z���`�r9��-�Q���噑"�.,����!�jyϴ�a*+M�O�'e��H�X~9�vՙ��sVd�4��T��.7��|���=N�Ux����!1���OӤ������3ς*����Ip
_�<�L]p{Ӯ�U�-�!�m�9���'g���Q��0x,L՝�`�d7��(ZD�Z�H�'�7�Ģ�0� A+��֌X�ӌ��M6[�W�蕐��Eӟ]�i�7�Yw��\1���{�Auf2��'�X��H�K�S.��)�j��Z��LS��L_`�R�pp�p(}=/�0뒡t���O�t�y��j6���qQ��׎4m%����7��Ŷ;�U�"�(}|4q��U4cw�x�#����~�Zr)�!�3��(�ec>V!�`%
�n��������фs�Y���߲C�&�
D����_�ג{!�.�[����T��Q6	H	��t�6y�8%�N��KG��0��_�ܰ�c��i����+J��*?Z�4>q���ר[k���{IJ8�]�0���*ω�_���Y5Z�)pGs&�3��l�TW϶�CA�Pg���(y�3Y��jz�K����-��*2<���m��*M�
�w%Z�(�$�T�>��@zBUɆ��Q/.�3 3%������^��Î����UdcU��� L/���dH8^�r~54U6�I�K%:C��}�g���
�_d�1-[�Mⅲ!L�>*��pw�F��S�oF_�8�Ğ�Dì؂��63�c�p��]�44&/���L���yYOD�Rm� -js�C�4��\N�5RO8q+y�ɘA/P��v�h�*��z�f`O���2�#:A�`��C=��μ*�VE�\���"!nQ9�J~��X���m��+��*Zeβ�׵c����m^����S�ɺ&�Ag%Cո��+�y��n*���b�q��,|Q�xB��rR���~���7I*4�ΎX�a�t�����i�V�R���fC}�za��3��f�����]��]��8��d 	�FpN��������x_f��!�.�TͱhA.�*����M[$&%�U,�����=�������f��@��or�=��61��e����2�;�I6�x��0Ǡ����%�syr�d��~	��z�D�� c��O���o=u��v�Ȫ{웃
����l����`�l� r@����9\zFzꆫ1�Ap���ϕ�e$���A/�yxP?�P��*u�z1%���f�!�i���-������.}-�+��)j0;��w��tmv�����C��ϴ�\�v�;�k�eS�g�+����ĩyk��|�k�%���P��G���-�Amp��]�I���α	��z�������Q����+s�7?�,��ziX3edQ!۷�s�g|Q_��~��� ���(��%�� \�U���&�K�x���$�,>,*��0n��M#����+XS�>>�B�j�����<z�5�3��bc�6zS��}���-
�t��+{�a��vγ�����ޕ�咢�뿂�%�F�'6�݂1���?N�ȴ�m0{v������X��G�Y�L�kR�r<��M*t�r������;uX�,(݇ٮ���U5la��]�PoUL����	�?FbuY���6�=E���q�u�g��+�R:^?��r�K�x.�\��֤5���ڿ�?ZJ�;���g�:>������q���yk�k���q�n��V1��������l`����]��F�;���Z?�$m�{��͍���c�Ew˖��b��m�%K��|%��J������-�à�����j���dOv�f�t�%��Z	U���&a��l�F^����:XR�hE�z�@V�@����8~��Z��X.�s��%<�e6������5����v������o�, O�M2ʪB4PZ�@�ñb�Ԁ
}V	��K��Ԛ������ve��M�B7^�0�(�/_E3W�[�q�u;�gT������3&uVi�'%t�x����Ќ�^�f�͓�֨���I����	tH�r���Zk١��no���8�/ТG� ]Dp�?��Pa�:1v� �z�6)ǀT"�`
\�+b�ގe��*D��U'濯R��x>G�)���<�i"�"�pm`@R�T�������*�-8�a{�i+���aimsG��z�4�O��+�Qn^8�Ί��b�{�!�<>ľ?ڏ���&AsF���v�(+#0��83a�lII�g��3~/�,���F<¸okm2,��\���t⬀{Z&���<q�U"�ݛ�"8��}l�Cg��+�����0���j=M����i2�F����_7�э%�WY!X��=��@.=�SMϴ�G9xl|����d�c�/�#�F� b�F�q��ʪs�8;�) 5?{
7���=�܅ ��`�ԧ���T�M/;�g�:�&	b;'3�Q�D~�w;���P�`��"l5�\�"��r�G�5�p���L�<�J����8��l>����E �0�$ү�W?�IV��tyꖇݨ�#>B��Õ�K�Vq����X�oE㋆OH�ԯ^��tl1���ad�s��K���nۮ%��R9�-�/�i�(�����K�S� �H���zq�ǪS���Sa���F�<�x�p [���9�y/��}���co��Ts]͡�����j�y�_5��OҮ�N,��`�w�QF��x#8�ȼT����ɬ��Նa�=	r�$}��uO�/6�VS������z�?D���G�~�aq���LbT�J~cP-pAA���ˣ^��P �ά�N����4��%�ݰOU�?.S�=�Q�W�B�����2��)�n0&k���:��ׯ�ɩ�5}���@��* �u�i�5(����0�gT��HN�4�}R�G]�"J-4O��/t����1Z�?)L�]�\�n�{0H"�͒��,�������z������:�'�ؠ"�.HD*,�=�|�r��6k�n�y��&�L\�P۬C��P��od
���v\�
���z�!�|�Q��M�X�2�bL�A	�@���QV�Q&�H�,�Q<벬"n"�:҅"O�8��[�pT2��l��Oh��'r�<�il��܎>	�^�Ԯ�˶oU�+`��a�^�#��T#��b����m}�t�,��2'��h(��2�jX͒�cܢ��(L�C6 ���0}[}�n���sY�Fc~��WK���c�j*���O^�ղp^�dwC$���-/����P�@�1�2��= �0��r�2\�\9L�� �Ҕ����`���Y��8`����D�B���\̣�+^���*4W�~O����>���O؈k&��g����C�U��0@�%��wr�F�Q�.!-��D <����xw��ߩ�Y�� �����Y�t��#�ΐ���.��\�P�!?�����P\�s=��Ry2�?f@��r����.;��π�3FR�&�pX:ޓd��3����-	�.�/I1��6����x�� ��9`�Au���ы�sx	/�#�g ��ޔ��jG0����60}\�W����ؑ�Hh�M~���"��>��}>���iy3��笀�b�=U�_`hM�mL�5�4�����k���$��	!?�� ����P�������n��[S�
�x�jce��}�7�Dƈ���7����"-�Ј��C��D;��K��:!`͂F�h���� �	C�6ta�⭍vT+;X&��"�d����W NƵ�*�A��]���V�YZa8σ�0.������M<����e!ۨ���ħ��#?�1�2���7.G��b��J�{I.ے�
%�B
6��O�O�@��殳��Q�ǒ��R��vn�p�ʄ�A��m������4߃^�L/�gn(��#���{:yI�8�����4��lg��V�$���޿iS��z$�ڰ�p��NJ������i��@2�+���0�Wc�;��%j�c��a��
جu��p�HZr��Ӽ*#�ї��
�?d��P�E&)֍��ȑ���,@ˢ��"�
Ͳ>���{��.O�,A��)^b \R�;�ǁ���5���� $)�v׆�I��о�1���E@���3��e$˘�=���)%��شL[�K7]�yo�CѼP��R�/�<n@R�;7χ�@��4��$#z||�B���<�0����9(��8���2yɞ�Q/���Ҷ"�yb�>��-�bF�f���Ӿ��&"��#M�7��1�����k	6&�����2L�i���7�X���%�c�wꖝ}�g��[�����P��zB�M`[P�Aڔ�<�z�(�S��H�ʒ�k��8`��;AW�ZZ��5�z]c\��ba�!��n;4#ܕ�d�_���.���T�l��H��Q��!%7��4�KM���Ti�(`C8����a�܀�x���ȢwB�]:l($d��YR<�;G�����1�:�w3o���R5�%iz륞1�%ە��<`�e��Ha.�3��8^���� �&��JAE5�ٳ�q��������5�y/}zZ�u>��?�K'��s�H����_���=%Xa�Ga�^�4�F�S���*��P��oa������D�i�r�NS��k�����d���p�1�'ɼ�qo[�^