XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����zу�45f�����N7�ɘe�Z�;?	">�M��Ľao�[T�W����"�+��^H7Z�
�b
?�S,yt54Y�Ig��S�aR[��q�*D������8�����ݐ�K��$���>m������[��e�����͊�R��`	'/�k�N]���;�G�?�3�ػM�C;�}�T�D@�ʠ�U�%�S[�'��KsE��yж�5ۊN@'��| ڀ� ���/}i�?��ϖ2� �������?=��D��O��D�Y�i�hŝ��D�if��`�S,�w J/��������#�Ƃw�]0�P!��X�qo׊U*B�!��=ɽ;��GF�#�T��n2����<�9o��Sy�ׂ�u�1�x��s5���|/�R���e��tj+��08�r2�5�$w[� \u�I�y?ۊ����~+�E@c�{V� ��Zr\<.XX��4ՈL�-AE�l�.d�wi��]��z[�}r
N�<#�����2�4�:׬d�`w�"֡Nz���/���Ӽep�K�����i�LqB�&<�R&Qf����G���4���R3���9ˢ^���wld	�ߣ��L�����P�	h�p�̎`sB�m_!q��d�n�/�0���8���-m�锺n�bm�����r�Yq[Z���ww�]��\�w�x�ن��F�y�+-<(����ć�t���D��J��!��|��j��o����)¸"'Im��?����=�H�ү����fP��t� z2 �z{t�<U���XlxVHYEB    39de    1170��I}Y���v��AGSE���kF{^p)qC���9'�X�"�>�T��H���̗#�PGWʻD��ܔ �(��I�:�����W����󓩋{S���JoosC6A�@I\tp>6Gv&rWn w-T���˛��kЀ��9��h�+������zq	?��L܍+��k�[ ������d�R�\�? �K4'M��|z��>.�}$C�_���>o������g��MUS����,(�.�X�Ynv�d�n>�PZ��Dob�a�"a���1{U�.R�M#ػ�(t�!�~{�A۩�o~��q��)���s/�0���/�,�m���|S�	��
���C��3���|W��"���z��p{���� [�D&铍"�hx��P�aX��-įHO&�����8���kf'�eFQs������y��5E�<��2{�[�N7�&ݾ$iSb��.냘�ࡻ^��)����]F�%������n�+a?#��{�C����S#�8&,N�i���ؗ.F�Q+�%c'��@����%�o%�Ж].��
����k}"�a����L�g����59��,�~�`�-��*��5��������GX�̉�NGVx}:.��7S-��k����a"n���P|���ء#��v�8���W�T�P��'d��|i��O�>���!��r��_��>��^�2I��('X���dC�94,K�`�������b?�xg\�8���ˌ]����A�2AVC��:�|ə$��E��r����;��qQ�V���E�.)l.�����Z��:���t�,�K뷌�}́�I�f�p�\@5��;ďK:��I�Ad'۬;/����3=b�}[��yhw��ʨ��+)o�T	@<��\���2��j'�2�G9?j��}����R.�ʦ�x4�`�cȨ��kV�j�5̰�F�����)���$[�U�`��.����wOb�T�/"�IO�u�J;�(��� ��c�&F�w9�����q��a�4�wߞ_oѥ?�><�"�n���)=���"(9����g��-�j�wuQ��W�Q�{�6�'�{s�D�7������sT�^6<Vr��'�i�b��@�����NI�e���3}� P�!���R��J�9�>���	���,�^�!s��]��Y"�d�8s�X�t��5`2p~:�L�-S�=1X����7�}g�PS��<����4g�ys��mԄ�52�ٳb3G�k�������'�h3���?�Y+���4�P�lz��&z�v�Ǿ��\�?E�m$���B��K��c���>n�}��Ia�����GV�����-Go6��[_�����wf�^�҄�ƒ�NL`�p��^��.���Æ�w���\NV�t����ݣ�ܚ������r.��E�2���gI�p��ĵo��	���J�B7�<�L�MD2�nH
��|��}[~(�xHʩū�8�3\D�)��[=�ҍ�P��{�пQt�L'Y��=���J��nHPp��O޻��
�;���L	R{&��B�}[s�PX�:a��BƟ�z�]�C�(I��a-�6?NK�� JI�����ө��P�͑����]���T�D�U�'9o�bz��<�����kY�q�i�g�o���m��0�"���C�T���'vϻ�o��d�����N�PH�a�c�ϊ���K����1������g�,Օ�-;�Ab�>�iz\�=c /&WWi�!ڪ�DU�49�wXšt�5g�H�%�"?j,��K���V{�<�4��~@�w�6Tg��dC�(T����8� W���%��O؄MZ�7�v��������Z6�d=S2��H�,��l�V��l�ט&�N~Bα����Q>��R,9�.H�l���
}�X��}y�R��#큯L���W�է��4�M�vkm�Sɚ�"�\5AMT,f�J���7��ܒ�t5�N������Xu��%(~����ܱ=�9�A��mlBc���T�|�h�{��f��p��3\a(�K��X���z�1)L��Y��r?-��N3_����#����5�U(��W�bU����\������|�!����f1Wt$T]	P�C�_�6s��o��C�qZ��tr��H@h���{ԭ�جi���|�%7�=����nw�d�k�	v��!.&,y$q�m�=�y<
[�#���AYUŨ.��ϋ��`�[M�R48qP��Nt4s�O�Ӄ��(H�5:��"?2���T���O+�]���d�D!�,�M5���Tݮ���"w���/�5���J�B���_�fT��F!��}m6�t�
y�A�� S�Y�������j����ǾUA��6\����.
6lBI��D�B�:�J>�v� ��6�M��n�+G0=pח׃��Za9�=S�
_����Ԫ��o���!x�a;�z'�i3c�'�� ��%:r�����U=���W��8F�y>G�C����Z���o��]:��2qj7�֮�m7�>�	��sG��)�Ӡ�cBIZ��zYU��T	��Bn���3F@�鴏|'a���I���΃7�=�����\�b'�	o��kQ���� �R�E�����L�n�:!YJ�>Irb���=e�Kq>���ԥ�)����" �"$d��#̐~*|��T�.
d�� m�� �Xq�j� P&4�^�s,.#k�Չ�%�9� �䋲&$8\�@�����ha2PIǷ����bʲ_M�����lJ�t���!�&|�]W@[�}NF\��rU�[�j���=�Ս��9R�2j�Y��/N�g��o�)Fe˅�� �4�(+�KH�l������L�@�	6Z��q�L���n��F@��i~��3
y���=�U{�"�O$�����I��~����o^|���ַ��D����H�,�8�U=x-�'�j�.j��/��{k�Z�x��2r��ǻ�T�hy��[P�����}a�y���9g�m_�}p~H|��=�)�Q��I����Ž{4Æ�����'�zD�m�o�:�~>���8z��خd�$����B���MI��l�.Ps�z",,���!���L4
BǼ_[`xhV)cn�d�鉃c��tÉ�H�Y�2`����m�x�U�|��M����J���L��zU3�e�u�
�~��er�n^�v�e�aM��˽v�����u�裶o��g���<�\{�#���n�5J�|�0F��؋�wrEl����>�
�t4S�96���?�"�#)X�0�Js$���O�G��K\���|� A�սk�Q��d3�a@	��TU�c&�n�j�;��`����Jj���7�59�<��T��MϽ��+��������&��3�w�B�N����@���M��c5ʽ���ɥe�/���M�4�S�Ӏ������k?��xhk��"4���e�B��!�=�	=N�F$�ş
)N}Z���ju%|�21Vќ�Gs77�������g��e2��CJF0K9i
W!�TC��c����W$"�Gn��ˆQ�)�S>�GUus1�ٍ(@�p2J��#��J�z��L���r'��x۴c���^`l�]�kǅ�PIL��(��\�3g��HS�lN����^4F9��?r�W:���c�M�߃n����成�`��?��� ��<��K�|��1�NQ ���Ԣ/� 	�z3$����j��MG��g�O�:�M��(����;�m��q��.�t������m�JiĜ��+5g"zW�ʐ'.�/@���@p�k=a�%ː���UP2��vk$Ͽ�09{0�F�O��"���k���o�[���:
��`~
!�|0��o�[����0+׵%��bB�&S�_'X�����>;��Aq6Q�O��|鐠�4 f�A�fe;�����})g�nf�Q���s	L7l>�xqhb:��VK�(���P���j��p
n�P906��e��5e��&���2~�&�1cr`�uz��E@P��ə�tR�qe�>���5���'zkx�������~@���	��4�n��ۻ�V5/��Mg#59Z�w�[	�F3J3}K��m�:�9�����0�w���%���ʹ0]�ϋ�S)���)��+m�a�[vy� {��M����<�y[��-�?��.-?e�I?��R��B�>3@Z�\4tkfZ7:F%v�73#����^���Dh���ܥ�aS[�A�N����^��bUL
ԦD:}j���o�	��t�G�f�h!��s*����P_Y3�^�p��4���wGB��Mu���k�1*�˦�@�n=)�9�`bH���
��~�=)��9i$[�G�
t_f��H�^G���������3���e��S���x�L٭:��