XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���9�鷀(0�a��뗤��]s����w�	_����Ǵe�?�G'FB�ɤ��tRBR4�O����-�L!�-*�(�7�5�ݬ��0Ӷ��?h���*��2(R���<bnf�a<̭����~�x���9�s�m�? R,�p���j�%�D�Zb���-ni�*�L��;~��w�_p�K���f��?N9�/X�\��7���S�L�c!Z+�m����6��bRy� �@�p�(T(�͞-5�F�	y����PR{0E^+u�B<�BU�9��l6=����س���q�U���/��ҝ�r<����Ʋߨ��ǒ��P|2�w ř\�����9��F��%�����#Z�z�=J�� �"��~�[�F�?�iy�O����x	��X 6-���cd��FP Vi�<4�|F�G��-��5�t�״��M���b)`|
]3��<����Fh|�s83�6�0�'���߉c�ry�]CU�#�KD ��pi�0$.@�$.0�c4��{�*6\ȹ��7�"��;dDhLա��۟:���r��M�����oaГ���|�`vM�����O��kpj"Ґt�d&�:�WB����� �o���ؑ�#����3�^X5/�˿[�V�U̶u� �j�vuG�-����}�r;��(E��A��7/�D�ش�Қ�tɱD���x�VTS2�2Z���6�r�(�}�Q
Z�&�o��n��-tX�P�>rwl�l ��es^�t 1���O�(]8��RXq��XlxVHYEB    374e     ea0�}�ٰ^(�Y�Y���^TWk#dT1E׃t�~:{�/>7���(��Mr��D`�W���tG��̕�G�[�u��g��3|.�%R�[<���n4&t���/�ʙ�:<�{�����^�K�B�P2�l�t/�BA��r3�meܰ�3P@��o%����U:H��Up�N���j�oХ��w��"�{����(A{ڟ�p=E>;�_��G3R�̇����v�l#�i�^��-��-V��9���L&�B���G,In�b�"�w@�]K��?�6�Z�T%*����9
J9!����2�yM|5��0 y�	��F��޾��C���"}�ۛ�%�P���R@:��)I�q�,E?�B�8!b���`|7�&,2*�?�;���[~����(j�����AM�(Ou��2[��
 ��Rm�#�{�t[~��Ǐ[��������쳐�z3����\˔���'r� ����'�Q�8��,ۃ�Tv�汘�$�2- � "{��@��{�A��D��
̙i�s�.���iC����h��6u����C�Q�?���!P~C���{ᕀ+I�u�3OmG�
ِ�ƾ��ː?�	D55B�R~��:7�d���Q��NwC��~ ~(6����pV��}���V�x���;�=��ǚFv�%;��@�z%���%U���Ͽ�y8���B���q1�[�Z����r�r΃��T���-O+/���V��9@��p@@K4�Q������ ��ϭ�@Xp��E.�$Q\�����U����)��a`b�CTe�ě����94[V��5}������=���'���\|c)�$p��EZO�o4JO8$�7,���~t~�f#,��+8+�Ƴ~H��=t)�خ1Zu�8�L�d7C�ǓKE�;�d���_�\#	��{7e_��>�X~�c���$)��O
�с�'����wD>R���H�捣_�#̘�3�&��n���0is���=� �m5��S\�6�8�a��wJ	�D��{^?��e 4Ļȵ�P�ӥ��v�wB]ӗDr��K�t���{�����!���S�K��}'�h>����|�q�}Z{A�����+��ָj�a��&��	-4�h;z�9� 5&�U������QwZ'�"� �f��=��W�}��:}��1���8W�`��F�D�恑�|�~��`X� 'o,�L��_��7� � �1����K��gՌ�Uu�,va��1��Y{��|q'�\���Y�S`fn}�7 cV�&<KMք[�@Re�9;)/Ż'*,���b&��X���S�������+ (�Zn�؋E�B)!vd����u|͗�ҁa>ۋ2�*�ޙҶ�%��, �'=�ý�Q��������ޘ���5
[ݙzFI1k���P�J�5��0�'�Hx���1C7���K�;	J���*�9~��^�V&�j�>�1|�5�-m#�'��(P��uXo�n����;��O-ɶ�*@�Z,�ҧ�o��oV�
ދ������9Ѷ�EP������(:n�[�t6/�l>�8#ӽ/G����'q�Mg�W���J�{O�T��ۍ��՘=
7i?�jN�1��Y_��Y�^/����d�u�oI � �ʰX2De�FO Wg"�zi.�F!��r%���߮f��h��~��T%.���K�M,��0)r�DL�[�;�����+A�����*����_s�%-�� s����I��ؙ�僷�U�� `7��v��>���l�D�¤n�J�;uW�j��c���#��8ō�m��y��L|2�TƘe�c�犳�P��������2+홋�"�b˨-�R&�>C_�pÕ�AF SY�ЙzM�>�+$u%��f)�?�y�{K��ݭ�[�
ўc-ᴗ)aE6ІZ�E��������ϬѰQ�d��[�Sy%��z���]H_qŴX�<����=����	+��=�Eß�^7I�g!�wb��
p*C�/�����u(D���������,�AW��;�-+P�]�ϗ��
9��f����kh#�O�51�O�o��~Gxy]@���#&�O-���c�hm(���qۄM,2CM�d��eۆ��x�<3I�ֱ���j2�r<�xdX��R�R���q�oar�b}���x�JX߳��mA��Fxt~U�^Y��z���q����.�M�G�@x�)~��v�go����`�2�E�;R��>����s�n�Q��; 8ߐ�~�����eJj��f�)\G~����̪�	�x�,|㮸��R�^�K!Uh9Z!�r3�gh��BC���S�x'�5I��v�$�q�R|D2T��]b�6����:��,��!��%{�r38���	7��Y�Y#��e�����'�c����>������#�r���a�A�MX�J$z���@�@��g�Oxɂ�1�-��􂘧]�z�6Cx�rT�K_�UN�jra��qq�I�o��u���M��>_g�̼��knq	+&w��4��?�Y�?��KH7�W|O���3݋?X��ﰖ��wT�����l�%��:%�`����I��A�������)7g��:�_vF�WF�)���훀����7nn,�	BD���gH��-z���qOV���e�ױL�pY:�W��խ��A$������*��9�m�;�)7�r�*o�zs�x�AӦ�h���4��J�ao~ܨ!�\5I3����`EX���P"_�g�$�;p�x�u�P>��#���`y��qr`X���g��Y��Y;Z���ֳe�|�d]��v{6ؤ~�$�����>��m������ݞ�>����i`Gk5�g��Vt��C�a�j<V`[X? �ůL�m%�������Tʓ�Q;��%����!A��D���sj>ЕN"�F1<`��#�G��ڣ�ǒw�|��8�O�k0=�MrX��I��߰Wc����-���+�
_���ag��	V��%��u�(����߽�b��x+��{ZD���B0�1�}��}�����i���.Ԃ� -/o@����
�	!R�\>r�`}��@�(c��ⴈt�JM$�;2�%�m1��t�I)\q����+�V�K:!=�� 4�k�4�?"8��� ��cg��WX����Fl�НS<TQ&o�w2L-��Qͪ	�)[> 0Q�I��
,k� �	��4+���c�ɨ���P{,�	�½Ѕ�f�m���@ި&-J���StDN��.��22�M*��@l"+@�q2U�.�􋽈�w/eL뒓��������� �sRL<]�Χ?�8�!�X%��]��m֖�,�.����#��Icl�!�amGg�+�i�s���w���18-��[�j��7aqZ��/�gȽ^rK���h��jS�Z�)�����4r��M��+k3"�B{0b���� 2gi��.A���_}�l����z
]汨W��9.�Y�G�=1��aqRzv;�g� �7���kl>���thx	D��RQ5j����q������%���\RB���_32~��eS���[��������jas�Yz�����L	e�&*GT"4ݸR��M��'$�r���*>[S���iɢ̶TE+!������\��ު��$�\6%\�'��ދ�K�#f��cA�M�Z薂�+Kȓ����H/]��b<P�"