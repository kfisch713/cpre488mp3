XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����ԉ�E[�6�bu�a�q[#B'���}�$�����H��&�|Y~�<;��/�9��vzY�������W,0(�B�H�]3L�Y�s�re�}NI���\��/�u%F�-��UcBlv�+Q�A��9�?��a��/+ʺ��vGf�b\�s��1b��E�ʖ�x;_;������\��3}�?-	o%o7��J���E[S�ݳ�t��v:cU��A
[x�)�f3}�� �~� 866�_<�{��>�R���f���D�����ŃwG	9��}�,���5S�!ډ�i�*�@�ܐIX����<eJ\��PE�~`u7��H4�6F���g>�٫�������R�fJ��y��H7�i��H>S�xD�aєR�ʀ�(�Zj�iLN�'N3��y�txO��=H��@��@�O0�+Y�	s�/�����ٽS#^첊d%8"���<-����G�~}�}+����kT��00���"6*���ֆ:[ղ�k��O��Ɵ��:��zw�b�af7V?��0�j��umTo�[�tö����ݮ�"�y�F��7����	��!��| ��&`C���ąj
O���W���}!�7��[oc~��|�m�&5�l��U�o1�;��y���$��{؂�RW���I�.���Bb�C��
�ጇS����yW˓Ҟ�?Ǟ���-6�������T2�	���$������q��$н�	�5����4�>��9�j/M����F��7>M���XlxVHYEB    af58    1ac0�@���:w|pIl!RT����F��>�e�9�SjΓW=Z��#����~S�b<M2�0�`���������R��*����F7����l�V�23,��!~����t9����viD:j8�q{;/�H��Cqd4�+[s�v�w�}j������˳�`����zp�lζ�J+=g�c�.�$1���羛��h��1�7#2��F�){�bb�1�A0M�M_
�*���囇Rk��t�2�ݏaZ�z_ ۮ4��ǡÖͨ�y� �N��J�;�� �R?%�wd�ɂ�M3&xw�"�IVoOa(jPWKg���x�h��J
��AD�˦�]������%{ϔ���=�����:�)���g��'1a��~><P/�sX-A�=��t��$�K�)�<�����5Z��:=�UU�!c�M#�gJ=��UM������WTqlk��T��8tJ`d$�8����3��c�W�'�+�D�D�G½ dK'{��NQ�x��V��;宩�/�+�J��d{��N�#H���Zg�a>陊�uʏ+�F�[#L	=�8Q/ƫ���C���m�E��!�����OZ���I�����9}�,��P��+(��)��g8���W������{	h����I�5��l?#��tjv+T!K�����]'+�ٸ>Ào'Ò��X�J�8�7�gv�/q2��DD��K����g*��$Z�Ԧ;x����D��v/���1?�M䗃GH�Ԥ1��6.�E����4��{mם�����~��#�\r~���ج�Ū�!�0+�����,���M���<�sU� |L�L�#vd&��.�6e��ε�҉*��q��xz�J
���T��`�:<�4�(G�F��]�W$�&������;sT{L��{���?�0)L�Fŧ��8}+ϩ�&�l�D��ʿ��j63���̼ni%'}�F��%�4�U��(�2�[e��v�D��'���
M3�r��:ՍT��_�R�^4ODٓ��K�(��#��F��Ӓ�)�<���� ��Ya|s�0�*КF��$:��V�g�߼�D����;EX�w���x�0Fn_.�A��s�H��'�� !0�޺�K������v��C����	�"DZ�7A�7�8���-oa�8���'�R���[d8)WR��3NųP�3�*�fS����$���` �n��ف>��@w�t��+�:��R��q����ej�[�Y���s�s���� ��_qR ��R�>��Ʈ�U7b����qR���ˤnA��n%� �u3#��\=9�I�t�˫�Q���j�i>ў�҈�#�喱�/��a?������d!x�͌�ۼp (�^�/H�Zɉ 9r�ka�j�URmσ-1[�d��DR~�C�"S$)l������{��C�8U� ��b?����-��pz�5N�t,&��OyV&"i)F�1����E���Ҽ8�O,�6{�5�8䊜4U�[��Zz��`xA�溤S���U]hq����#}6.l�=�(q�Ԍ���#f,:�}�;u��׾׿&<�?mb1C�%���ERr�ϼM��44yn��p6�Ҿ7
h�Ҽ@BD�n�i��N�S��;F��R�46��1J��L��f?pIp�h�a:2d�Z��hD��_�j!E�)���Y��Z3.�
��ю�	���NU	C%�663W0�L��neJ�'�ǽ�'��w��H��S��o$ğ����$Z$�ه5��o�4f��|M&Q�*3XJ� �8����W*� ,�?�&,{͗��Dw-(~�RY�0������0������E����r&�g��k�ߍ{f�g|�@
{���>�6�Y�`b��z�Vr�~�)�U���	��.:�c�3���
O0A�Y��N�-D����ǜ��c1!�u���p5h��b��u{w൘w@�܊�l�#�L�S)���q�����6y��v����(���x��f$��0�[���A��j��&uly�܃C��)5�YN�0T	�Dw�Fe>�] �|lU���E�J��N&���L�l�6Ho�(�r�1�
li4��y��$�������6M�^ܼ_��=ae�C;���e��RG�*� e�����W��/���>��*ES���L�VYɈ���q2L���s��{@�}�����6��\t},���0����q*���3�q��_��-�>FS��h8���e���bK��=����A[�ׇ�ea�yE���M����O�w۩��#�
��.A�S8��>��~���fT�Y��+E�b{�����q�l�NH�����g�W�ܓF�w&��t����j8�Rsax����0���jW 8j��IX��c�GK�*}������X,=�lcJ�1^�#
�S��g�Ч� Y{$x���Y�x7��h�d�jc��e�-	""]w;��2��n���ӹ���~���4�@�S"�����>���%p�E�/Ŝ���	<�',F��x�$���X��u�&�\�қ9�(}kȒ�꿦.���A����@�t5��XӃ�ւ�鯭T��x$�(��,�TB^������ R��ko�
��'�`˛e��QCA|��-�nnT�L�}���o�)��Z@��E�F=D�<�+��iR�/�q����S�s�F�;�g,hBM¤h8 kX�!��[k?i���Dɺ��U�#L���V�j$>�X�ȼ�l4��d�ė�:$���NF�q�Wxcx~��kzM��-���!��8�Ԁ���N��2��3S,��q���b��0�|B��\wvƽ����Em���	N4�)���@��Z6�z�(�1ߺ��o�/@�C��:��;�U�`-;�Z|xT~˹ʜ��=���ڔM5<��i�����/�(�yQ�)����.	i�]_l*�7��b����v��m���F��{��!,�]%u2�/C�zPJ[�5A]C�*i�����y �#*`�s1]�_�3V#��5])�9��� ��E���S�'��q��J�q��Z}�������õ�Z��$��j�G	�ף�����vM��kK>��@��L�TE��a<Ƞ��l�Kgȴ��HY���q���.(��׼t��״Kt��v�mؖ�c�a����P��e>��%M��|	Y�v�C�I���K�	�-JA�y��%�K�a����F�'dW��t"�䰽&.�����o鲏��k����i�O�S����˺��c�zt�`EiƠ@��M拝�Y�v�/����a�RC�3.�N9x8Ts��֦�ib�����<w���0�z�@ՁĞx��4�$�"*��m)�٭?b���}��|�JN��N�f�lnǝ��i1 Np�H`�yͅ�����H�����)y�zJH= %%�!ƙ%�g��K�>6�� ��ُ���z��͒��M4㸲�_�+��#{B�B�����ǸX�D짴tsay8����e!���raj�'�ȱ���S4;��폣p:�{t'сq^);��D�v�}�۝�aU��Q��!�[;��G'��yZW�!�M��@�Y���wvB�O��&�}�z�L�Z��HӘ�A�{
U)`���c¨b[5��}l��O
]`�|�z�6�7�[�����fjK���{q����Y�#',ʋٯ;4I��Ӑ԰ҥ�X?��%%�<r$��$���Lݺ	�� �k�=wvM��*���OY�vf�B��~�,T���<^��Yǜ-_*�L�d�/Rw�e�%�u���2,D��O.��˅�iQ���e�W&�p�ez���e4sV'�%�,�_W+vIj`�|O8\�����g�8�~�tybklkВ���(e���yc-��vm��uP*�3μ��qOvW���U�8�+�:�[�Ѱaq�݊���/�-��c�S12w��Ul����n3�>�9���R����Z%��F��ʋ��]ä�Z�ق��J���&�җC����,�+���n7�0�q����p���6��`�Џ��[�c������
6}]�W����\�7�ΆYnr�[�!��ц�Nke��u4�|/����/�ח�E���&�X'
�D�Xgr�Llo�1�Z*xD�[�q/u��c�K�A^2��G2Gxٿh���6*�eVH�j�f"z�)+�:�J����v4_�]����.�4ǃ�)v��! n3�2�tZ?mxQ��@��Zp�n�Z�$�ٛ�k��1���C0aW��)8:��@pL�.� �I1�Q��l�pir#~����O��_��b��(v�T�����<��#��ڤ���GY�8�g�Dh
DՏ��aD}����{I��������	8Vw�o�Fq�ÚL��e���y��zL�Z�Ƅي@h%tR'Y�[/, �8�4:�Q��P����eE�J�����V	zw~VS%ex.��Y��'���/�����1�j��#���=)�u�K�\�����}��W�Ah'�v����fG�y:TO��AS�2i��?��p�W�V�qV��Fޝ�-*���c<�T
��sltI9xfߎ�uvk��wݮ��H��n�W�NxSe����.�7/u�{Ug�+\a��@
.x�Б
"�x���y	����l��t�9��s��糅�����$^�	*Ręи����s��DƎ�+_��3`'��(�͇Y�NSͽh͖���9�@��2��V���J_F��Zs�HC��e8إ��?�����)��{ ׻;J���.P��J��J�	���Q=�@{l%����>��WJ��!�����$�IA�.3��T�o0Rc�
���I
��_���;�3澺q�t�o����4�1<�cK�Z���� b�U�[�z���@		�BEފ	�NV�١�M�9}Fa7/��G(x��n�����	-�ů7V��H��VQ!������@G	^�z�K�;���N���\r�C`7l��������Pc:�£�"vh*0���h=�D!��"����E���d��]��gw�q�5pl�W��Gp�Hw=���7Sj�'c��0vʕ��/tfܯ���Y�Z��a�.ᴮ�$�m�j@�s�� UXs]�3!`�e�K�zXm R}"� |�¸Nn��C�LqP]�-}��,Il+�*�C�g곾tUf ���Ж��>4M�m�}�T]h��B�2��W�)^"��W5p����t���q�{��-���>=gj2V����./6�>���/,��=3��g��>�`��.�����MO�әHE,�;oܹl������j �C�D�pL x����]0�"��͡�4��7��J2I�F��+��iXl����b�7Ҥ��aꅛ����'�*֓�2��~�X�!;e"�RoC;��]h��,�6r�`T��+��_���M���ٿ�N3��[��j��y�*��{�F�.�x���i��JR��&����V�<,�F<�I��6rrO�c�؁7����ָ�㦕i�40n0�^�DvqG G�J�gE�*d0���y��=3����F�)���k�D�2ԴV�Tx��Q=.����s��UƑ_ܻ����^��Pj�\��Vp�D!^!�/t_FZz����_��Z]�EA��"�ܟ����;����C�7R�������٪��`:?�_�nZ7���W���[0�fy��뻱����g��.��KPY����~ �����^�厷4��t�U�e�d����=�ܜ���hO5���/��'��J__SZ*=w�qx�aM�Dk3O����=ip� _�U��Rm�	�|��@e������7��Xк'�F������Fy���?S+�K�D`U;	�N0`���Ð����/4��86���IOf_T��Z#Ѝ��T���I7p�đZK댈BX�(t�X�MI#�\u+j,���$1,�bpl:3:Yڜѿt8��S�Q�)����?��ܭ�%
.�.׶���æ2Y7Hv.��	���6q�ǈ�T�÷]������ܺ�`�*�b��g�M\�q�Y��UG�����\������yO.��0��~��iL�%� �.;��2������z�g�WU_KA)a��cU0ؠ�/8���z���x��C䷯_�^�� �7��|>	������=�BΠ�\�D#H��7�P��r2�PvXT�^S}�Ԕ��f	�sZ*��id������ќɥO�xV�.��Ђ{ĝ�Q��_"�$�Y��Q�ߺ�V�yԡ���t2���yp}A� ��_��՗���+�(7s�.k#B�l�@��k���S�}�/tj2�l���JU�1҃��.K��"����ax�����3
��Cժnkp��pI&�R���4��+)��M�<NFt}����6w�Ԭv���[��#_�6��]�=����.#����c�o���!H��[�^s�;��yN_A�۵�>,��T�K@�8!�7�K�Ⱥ��-����2��7���2�w��Է��`Q<�-��� 	(n�7�!��<N�Bzt�{�3�p��U
Y4�q��~"�Y�`�D�Q�k����E���da>���^���ψ�Lp�«|�R|啔���)JZ�j�&q�B���^�Mg��EA�������f�B���[9֊�`���x�YqkΆ��=�?"���k���Z�b�n�˺#�δ4 E�vE��'���v��w�/c뜸5����S֝����V�!���>��j(" ���tOG�/�E_�r�_[9hY5�|���m3��|6M��(c��u������Np��c%7�#%��/,V�#g���r"�}	��