XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��0��y3�?��(3O��-�����m�ºgh� �w߀Ѡ��Hgǯ>�<���H��y�L�\	JǩĘ~�~R�Ġ���&of���K�V2�l��{�f�ڹ���Sy��[ν&h�� -ݦ���KV��M�������c$k%�d���8@���N*��t�"A}��#ɻB�����T����&���Z���Ŷ�Mى�'����yX�5|Ɇ�+�7�� z�����͏Io��	����������+�/�v��;�7p���>L9�}�|�bL(<�חj�*��ꪪ�46t�%��}lO�3PԚ�Z�Z�e[����*z�Oe����н8 ���2��ǝ^46�"��0Z��їk�+�_�</r��
%{�U�K�o,��Hb�������k����+߽g�
uɞ�(��uj*Z�?�:J��t=?/��\ZΕ�۵�%$\��h�Q��oX�����-'Q���ً�\��ٿ)?����N)�F:���q|�x�̸�-�t����q7��2��4�>%�b��٬"�B	��Z�1,���~T���/����'��&�k�Vo�5�[��^���(��}�y@���Z�ǩh������ �|��в��Q�x��u�����7���
�!�����;��aB1�z;y��3�ŀ>R��r�^����A�����8��H��
�
Ód����͔lb�7���Ρ����ܤw\��W�G"�W$aT�
�A	b��}M��)��YJf�n��!#�7�68�"�yw�#,�XlxVHYEB    893b    1e30͒�\�K���#A��j� 
�b>pI�S��Nӿ��K�O��{�ꗮ>i6`��p4��r���s:���8�x��BG�9��<�C��g����2�%�oܚQ=���7|���f���"4���K�/p����U07A�kyq�p_ՁR�̡��k��U����:� V7V���)��]f`����xRܹ��]kha_����e{��'<9�#��>�F���%o�%0pv��_���E���I �ӄJ����tX��[x��\�J�fgc�q�}�T$K�W�"a�8[LI^)�J%-&��v�_XAE�k�eV�pX3g��3NG�{��q[v�ʄ��Wx$�mMܢ�'��P��˙y.��!���"i;u�:<e���ԥ�9J�#�x{�ϒ��wv����r#l����+�Q�)�i���D�7�n� `d��{��q���Զ�r�M�Tx�z��c����y[K3B��ݽ�Ŀ���*�;)�('}��!��~����:�h��:��6���6�q:���𕆧k�v�=�(�A��Ha����r�46j$ɰQ"}V����	Oyn1��8�p�����/��c�;n�����HD��H�$b�i�c�شs"3R���S��3}��]C�,�'�{�P�ۚ#��P�A߅�C�cy�E������b��~�7��`�<uE`m6�@�����!V��j��"���m�� ������-Wi)�T��3P�[��B�����)S�դ�]3����w���r���!�j�Ŵ�m��K����b�;H�>H���`�u�M� ��ɲf�2�Ꮪ'RG�q<��!V)k�/��Ws��#�8u�A��ټ{$^��2aQ�%� \�b�e@22��>$\:�{o���ƞ�:sƟ�k"��a/D�W_�hު�d�Τ���=4�Q���;�PR,	�*�3GLه��mp 4�>eX� nh>L�P`a�j�A��T��t�����\v�<Y�Yk~�K,W����b��0��I� ��3��'T��xjUm�5<0�xL��*1�V"ͨm�z�x)�Y )�]���Ee��A��&aF�/@��ZBa@�Ȣ�C:k����y^`G��+Zqg�zm�-��jH�"��(�ǫ����і{����� ��/�t���ui�����V0��&�P�8�S�ّ���ͽ;p��W0���d�U3Hm�@U՝���(��V.��)6��1H�M�$Fshr��@ˆ��Ͷ���E6�?9�T�G���=��L���-�r ����9!d`�~��db��+	���T�r����xV5oX���-�OKB�!o)�nל�7��}���g��Ux3l(.�}�Y��}�'�}�T!��bG�CM�Hv�����!Ǩz'aAQ74�y��n00�J�@�OY�켒.	��mqؒL��ᜋF��0@W���q?|���z?α������M0  ��k���y5X�b_��뢅o��F��w�
�c��z<��o;�Ƒ찇prt��ϧZh�zߥ��zN)�PF�r�Ÿ�2��Y�g�<#)O(#��j�B/A'����T�s+V��69���!��ޭ}��8�Q�����8�kO��p�)1S����k2/��6���<��-�����EX������ʩB��Ww6�p����>Yh���߿�s��Q���=h�^�=k$o	,m:���o����e3������t}DC����y�] ��f��a��Řۭ��h�Q��l@aO6'ơ��D8.�j������t��<� �ݦ���v�Ľ�� �����&�����]*��%Uoe�#a�� �L� ��saͰ����D�/ڊ�U��3���I��`��A�^Nn���R}����%lch��S���N�\�>�����F��'��O��g�U��I/qrz���Մ���R�����1EH��8�.h='�C���wHy&a�K���h}vg�G�g�6=L��e�xn�D�sgO����5OLI�0��mV��|��Xz�'�:��u�;٩w���S��'��K}�ɘ{�Ue��֋���I��2�j�uz{�X-�zHq°;�6�
hIN뉯[�C��6�u�NF�]j����{��O%�ׄ�.����w����$rjs�V���?�j� i+]�%4 p��aqƭ�4+���ɯˡ�o�e�|q���� ���7L�:��������m�h�����,�	=��-�l3fE�ܥz���œ�
��g����iȃ�-�50x`�qSX��|u$o��YK|;����Ə����X���Y�Ǿ,8KX��Ӛ�<���~��2kx:3�"}l��r[��_J�+ru�G����X��oJ�d+R�������H��1:�&E��.H�������,L����YXm�1=W�Hj�$\�����s���z��� 8d�P�?r�o��ޏ$��x�w����Lr^����a ��L3ژ���cy��2��ۡ�P��H�I ؍�m^:�l,'ZJT�1��Yc퓦'};����*4IqW.�&�Ǡ���(T�i�ݥ��*���:�X�0���c��Ь�W�6��~;)���A�G�T�T�4�h��9�tu��Ք���L7�+L3}����t�/�R�M钮t��6b�f&�7�[�n�^��UV\���O���ֺ�_�nC��n�zX�ɟ����|n	4v�/O/��w�ΤEOO��Ķ�ö鑎R'B����O�R�:��c9��U��"�PL�C�o��9��rDo���4��3���W��7���H��΁n�$�-�C�#f<<]�k"�ϻ뀎`u>�;�����E���D
��4�%8"�CN~�U��gR)O/��iL¢%[��O��}!��G	��j�l���.8�������òr8BVoR�[�U���	C"��qg-� s�)~��+1�><"���$m���x|*B�m<��j�&�N��3Ʈ����E^i��"��>�-NC
n���U뱘x��;^ձ����/�a��&+&���d���>�=u.?���s�ZW�\��[4,O<�!%Q��2��WW^~�ι�.Q�1m��zH��8m���CҤ!�p9�|���������Z0��m�@��rŞ+ \�����(�y=3&ENu"C�w� �D��LT�jQ���T-�ɰ��8��1-%�@v*1?"|�g�(�;-�k3_/Rg���+��2C��z� ��Ѳ0[�X����I)?�:��q�fsj�%���f۳ٮB���jZ��Պl�k0�z���	h7q��O�Q�o��D��܅������ �|�,���s�A6�Z/e 0�qaT��X��#	f�R��zUJ���F�����D�*6V��U>�,\��D�umM�N����J�0�m����uE;&���� ��,��S9/]Ј������)� ���(
Ԃ�RrY9��$��,�N�tG��i��>��_��h� �ƿ�Ć��t_3��Y5~O
}�!�J����S���{��[�q�5y�*�i'r.9m��5�##�I�'���w�r^d�W�#�^�>}}��j5#��C���n�6��Kl-�@Z�G-5.����-1�f�-�?�8/L��gv��������(EIBn��e�!�2�gZ��[�!�[0%���O:/�����.#{�+��a_�����(�뇷s�i�ch��&�0h��G�m�a�Q��5�gg�H�:��ص�i��j&/�_���qF��W��0���,{K�t�0�.��l�Ї���\Oط�{�!�����k�qFҳ��$�(�KZ�;����f�ˇ�80��5��C'���t�T��o~����K���e_=��%�*xܐ�r�j� ��/H�W���������q\(N��KUޕe��� �ǒ��BB ��5 Zp�#�E���t,߉m�l�ܽ�ȫ����`o�s2C*�eʊ���	�@�:�,SJ�� ���ت.���'��Q6�7�Oh�@l{�β~�3;s�$t%N���>L�t>�+k��1q��CJ��-:	�q<ŉ�����Ҫn��Hh�Z�I.�3���T�[���n㣵Y�J'D,�S���G��+���geɲ��:g{�A5�S:12F,=��ϱ�#���&�0�~�6[5��A�+��O��W$��M_��J[nΦp�+���,��|�(�C�۲��ϲ���O�iW�;������ɼysD;Gf^iVD�Ϋ��}�������)8�h�t��}�A`����6W���a �-m'��%Vjw&��1N�Q�D8�s��Ξ�\Ԇt�l�瀡����<7��쐀O�����n5�\�h,`�G�4s}��x ���/�A=���Gf"iRV�瓛����j��U�����m���ads ���?\_��BZEr��Je&�O�c�P��lOr�0&��Tih�}
8�*~�;(.�^��%	��
����]�5Kt��S��)leTz���D��~�P�g�Ư>c�lX���{X<޻�����Ɓ�t�^Zx"_��G�h�厈J!�%�Jۼ9��_��.�_��ʣ*k��A=l��U�U,4t0�H�^ʫ� "Уg<�0x�p���J�_y�����9�ڤ�4��	ݤ�MB��VdW�Ѕt�����.D�c�Z�"$��M/a7���YXӼs
���'To��T�=�cC���ub��kc��H Q�Ǔ�<�.C��\c�!pv@J��r�w 9�Z����GB�I�&K1�������ь�O�tcs�v��)5�sĝw�|������`�}��RA�<��Ngء����1L�2q���E��u�w�/5��l��<�s�����A
�l�N��m���w���qC��Vҝ3ZI�RٮRע�F���!�FfłJ�=e�xPv����p���.���,ߴ���b��Ѹ	�{��M�M�o���V��> ^���d�U��^��a��<�Rހ��\�	�y��%���N�I&�ɯ���%b�`��x؈�`#�t&�ϰX�0�X�g\�^���ڽ*�3�b��o2?ߣ޷Z��A����H��õ�s�h��ݴ�-9��k��ʚ��;��1_�� ,ʎ���D�Nr�U�!`Q�y��ր'J���#�c�x����#�A�NbJ�U�������p�4����@�Qq4)>h��)�mĸ	q�^3m����15{q�����3����]����M'xo:�G�}�s���PV�5���\2�!�v�	]�׼��Y%�$u��`�>`�V�9aP	M�o-.x�
�E���Y�Q`A�d�t.p��XO��§�5��_5/���!�=�qn�v1���MҰ�_i6&����	���(�ԆJ$N=�)��&����"B]�� ��z%v˕�ԯђ+7�O#\��xq��
�ۧ���*H��p�HrC�Q�@W��G��"G���~1JhLO�B�:���c��H[(�����"0��@��L��휿ۇ�=M%���:�(��T�J��oy������V�X��dˉ��I��U��t�Ds�E�Q�˥�H,��Z$Rư܍�۝o�u��-D_�4��fA�����/��,ֵU�����J�N���/��<��;<:�m1�>�M��9ã��n!m�!��e0/07��\��MK��6翕7I�ӍJ���>� rg����.�߽(�L���(G=w9`��i�?h�]�G��<�J����o����p@��=�.��b�.��K,�	g����lJ�V�X�
��T�6dgd�5��y�2f��W��{	�S,����ĳ���#��㭁�Uc�y�������#�OJ��.�
u-�3cS�AW��e��)�F$m5�:I�Lз&OO�ʉP�4���,v!D"|%)$2��`O�Ŝ�ƾDm���>ᅨ겔G�DJ����Jws{/�B.\A�~w�0P ]I.�5{��U��ju-��)���:B��ߖa�g2YX���7�M�,�3`oXw�T�Zq��s� =aph��^ @%lj�z�i��A�ރݠ�»h��MM!�e��¼����VM�S����,�����4A�p��
Ȩ���(���a�|K�8L�J�u*m��M8M@	�)�ɓf!�	�0kV��a��3�m�V<lʖ񯺑Pg��5��Бn�~j�Yߐ����σ��B���g�_`��4C��w�Pw� Q�i�{Ä$oi�9H����"dwu��DP��rgze 	[�|Z�kI�'"Œ%���H�O��=�1ȼ�$N��B,�x�S�/ �l֌��@ǲؾ�>�9��,��:���@��(�I?*��tlbSph�:m������[Ֆb*�Ls`�a�"��ɇƐ_���dʙ��d��CBY��/>�Wo�?|s��񐓤^ܞ�����C{�l�p�F������'��`'~�n�Sõ<\����7�m2J�<U.8�����m!4�>N0g�:�J�V��{ݟ�:��j%g���m�G��Q]c���s���W���.�0b��RI�t�t��4-�"o_FHWTp� �/T��ס�J�g%�h>I¿�I`S�e���&�r�<Cq�t���ω � �jn�g?��8
V#�c�t�zf�!�_^�T`�����%����A-%�Q���yo&h ?�m��a���Q&��N�!�s����<pmrC��3���8+�8kvt�8t4;�<�r&�a&�/�&���������7�й"~E0
hթ�!�C��u��%O��J�<��4z|��.�k����2�K\���Y��}�,
Y�,e#@��v\�Y�96Gm�����b��k�Չ}�]�gt�t�h�.4&�;��W>gq��p�lo�����B)M�@pH�r�D4u`���D���!�JG/����fB�BDE�\��zo&w�Rh>�p�#:i�4�0��� @��1�C��kabf�K��e�&�o����%y�!&ǂ���4��:���W:���-7���@��S�I��\*�|���i�U�(B�1e��6yB$Sn�}']bi^�RE����i>��Y�O�
fPƟ�"�}��XCN	%{��� �P(��儖�G:|"��`�Y��+��YR8��y[{���Y�/�=�O7�,T�h���/%#���Ш����g�6c��_���<�Va_��ɻl�c����5�~G�>C+6Z�I��m�2准�5��Y������	U������*�wm	5��[���-�T,!3��[t�\�}�<J�%��P�W�=
g2��T%�?��л�?�E���=M��B�ԚQY�W��Ǯfݖa�$D����+����s�(
�'M����_�Ѝn�8�ک�U���W����q��A��x�o�p�ݮ+9B�c�+�B
m���y�6_�1w(I���n-��#(��^;'��㿚�\�{o	<O�B%ǖNQ�l��o��@~R����"	Б+�<y܂�$�ퟪT�x����51��㺓�>��s�d��~\"(�"ν�V��w��0�u��� �����9H��r|{�A[��ڠr�XǇ�ҩv_��
�< �('\��&�$0�ݼ�z�N2~�.�Ӡ`x���z�,y� ���!$_