XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���]5N����+сY$��=�U�N��&7@uݶ���L�#L)q7	J���,��mC��vi�a���ٞ116tCw�?h�@���F�a�Sz�S#"��xN��ď2��k"�Χ0e�b���7�
G�P�q���$G��l@�z-;T������ʊЂ�T���NwW�{E�1������$�F	]�k4]9S��@=֮��-Rt�KK�i�Pb�Y'b�)�Sm��u�dE���(��@�'(�`�x8KP���
Ą��̙�)sG,C`F�l>���Ō��3YD� ����|�H�5���cv����Q ��#���'�z+��8���H4���Nz/e�^4#��b~�9�Z-�fHϺ��u�!+��.�Ԁ���#m�S�,P�A�[k��� "�����xs�3�y�-����~�XH�7�,ӑ�Q'%+7M���O�N(��0t�K�_�i��B�"��G�c��<��`����9��a�P��MN�O����a������u���P�Fq�/�q�ô޽�]��m�p��R����pAҽ�ˑ��L��C ���?2cY�&w,�6��)��ie\��E'2��.Eb���Ċ������_���2�I�-�zy�m���9�Ȃ8K�1�{�	oArͼI���/��X(�	{"D�L\��r9�s�J)s����uE=s�@¢�!�{�H�ZH���Cl7���r�6LT���_[���)�D����Z�7�!P\�Ck[�[���6DUN7ߗhd�XlxVHYEB     e07     680E�"�y�4<g��qb�Yg�S��uV���Y�x'6���-b�~X�T��h
`+���S���ɸ0��e���&}���7U�=��ޖ���'��X��؞~E�k~G��lw�Жuz����W�;D71��3���~����X������d��4�+���?S/Eg��
�?�x�L��;�Lu4	���e�֭n�_��O����%�@���М �����;k�x3 ����j=��O�'l�.�i�X�4���UW�J)��L��.�����	;��u���]��E��z7���}21�����$"
���3�o�
��w�����%A�P)���81;��G�������?9�z�|�-Ow���G�I�P�7�:UTF�����uJ��C�	����N6��L���%vK����E��б��c|I�P��[���$����fsy������J2Axi.�1�b��ۨ%�Fa�HB�`)���G��9 &yٺ�@~�J��~��V�g+����`��*b�N}Ll�Y�Y����4���$���0β9�q;�&k��2 ����.�VHt�H�[��j��?���_>l>�q��~��VO��g�6��'|�4`|�����1��=\�?���%&Cτ�� ��-5���p�ِ�:���L����(�������UW�LN9�����
~Lo@i�M֡񹧈�?*7i;��l���`�$N[�E����65k�������pǉ<0�zp����8���ϊǝ%2�����R_�����/��y�B��P�IlC|1�O`�L&3��zARb�Ր� /�]�!��a�k�:�����;0Xm�n�D�ȋ�O���4ۃ�����vt��ΞHTd��<�	{����?����o0��\P��Kz٠H��qY��m}3��R�]/k|�T��{s�Q_���A�#�����-��q�dB̉	��ޓ�(6D7c��o�ڧ�w\���!��?��&���*��fi|s��5&[��{VI�~S��+b���ќ��"��M��Q5W���$r�����֙+Y��@]��^@���S��J�(�w�ʟ�ݰ����#��=nԲ`iy�ƞھֺ�p�����zb���1+dǡQ�39��m�v�m
�ܵ[�F�,�� ���?�O� ������� ����M�=�>k�#�R+#�^N��e7�]��x����)�I�bg�-�5@���hW�/�d��W��b�� h����<x9�*|���ux��|��۵�
G��|�����\�d:����}��G��(t�S
�������z}ob�}J3� c@��l�;o���E���Y����G4��Tfk4��vf5���m\C'R�Oof�Qԧ?���YM�~ByA�
,J|v�Q�b9����2[���wr�9�M���4�LU b�E�W��0����}�=
I5k�2g0a�?"�Lmͼ�Zp�g���E�,a�uiZ@W� 7���E�W��is���r@Y�7��I�-/R���M�����0�c��<�x|�Vy��X7����ۮa�*8n�mTO�-�(�@��K�ξ���4
�^{֫��|��9z�C��T�B���,�@=�Ju4�F��(��#�,���Ư�!�S��B�N�+���K؊����