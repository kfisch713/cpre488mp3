XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����f��j�w�N�C�&�,��+J�E�=l��K������Hw�Z��*A�xzG�˜����n�(�]�A���*�,{�碉����6��Jd���IvQ��&�v/P�9c'�׮}?-��)��y�!s`AI����J+�ꁟ}I�v� }�n�s����6x��}�.�)�Fs����X�g��;���5������ٲ�+!d�<J�ZX̉\c�Ro�۪�|�,�]�p���g�`N}>F��"S:/�z��E߮#%0J�8���6_h��n���Ӊ�Tۤ~�į�0�"��0�g��������꺡�p(C�ݍ?^V�š�C����q�`=g��\��Z�q��F:vNد�U�N��4�P�9H�[�;t�;fu��'��K�3�3i��@l��}����}d�5��_���iuZ�w���򦇏}�a��Փ�������56���?�jU�;�E���aN��y�P�z�k~�p�NU�7��$�R)�����J�G���]��ʦ�x&�U��ȭ�gy/z�2���N�0&��H�呟���̈�]�Dľ$�YP��h�N��MQc��"���aԓ}�.�}?b�*��
p����ˡ��)�-�j�:h�ڑ��r�>����gA�����&�!	��];�Uْ��]�(�s��!�z$���-\��g]�
�;�ӛ_�]���֌�=!���ݚ(��f+��� &F�	��U$���V�뎟�=C`&}�Jv=XlxVHYEB    925c    1a60�������O�����X���H�=����>ī,�#�l�ؕ��F��q���t`�_�`�kN��{56)�'��pa�ϖ�ǡ��e.��d��(���ɑ�I~�uk�c�[�*bM��I�cܱW� l���j'�ƥ�l�>�.%���M�
M GM*�=�|E\J�"4���H�_�|J
]�R�O�����f�5��;�	�;�����i6<|���m��]�u�m\+{�*4�]��-D
 ���vK�A�� ,:'0�pSۼ�kxR��
S�&{�i�����@3e������m������٤༗U����H��6�������R���/j���8����jmUT�X!P|(�� !+���)Ĺ@aŕ���y���4��8���_�0�v�((^㞏ݛ6UC�;+Q�A��E����Xd�]$c�^^Hj���KB25�X?�*%�G�z��j�d�BzӃ~�E����;I8�R���?7T��X���N�2�~���@�+R�U�9�Z��Kw9����c>&��Yh�d8KK��r��>EVy���a���4w�*�-�s�4%��c=�;m+�[�� �Ƅ&q�xɫ��6���� �0鈊��7�^�?'�W*<���+	§�3>
�q��Q�*�؏�k��o�)[>7��.(�ye,��aN[�4�����0R��qƮ���"�G�c+f@,ڀ���h���B�:��)To^E"�dJ�cA#�i$� �1
� Ñ�-0_��R��V�&
��쾲Z=;�ɂcc%��I�����/k���K�+�����j�T�C:� ��\帠�W>�;߸��z��7$o!W"6Ö
��M�6�� l(�HרV�p+N"O0�s`ѽ� �	��ҷԋRF'_�ZJ�_S+RHeZ	�b��@yѷ/0��ˈ��}�����<��� ���O�)C�%��W�B��j��P8���; Ez��a� 6M_�ѐ�� Y	��w��x�H�raI��:���	��lk@?a����,y��*6U��K��'UfvK�`����P:�0��_�kq�d=�旳ܱ�*��՞��l<�.��˱�^>o����x£ag�iH@O�F�{09x�,��"Ij�����	@u}vuTS�Lp�{ӳ�!pN���h�N�h�B'�tj9Pr�n�m9��[���J�Tː�yr� ��W��6u+_�&5�#��w���������/��9�p�-�0Al���� B���g7�t��Y��[����~�������d��hߕ���ә��'3P�V���]�,�C��?�Q�t���Ѵ+��{�<��hW�\%Ni	��`�Qa&˟���C_97AK�n���"�16@�a��JA�𓹪��-��`�f�����&��w��}��_��P����]V�K��eL�?#$t�Qv1��q�'WMF?��bW�+���$�3�H��2;����w�>H��n]{"�xȷ�D���$�.�W�f�I-V�@x�E�ќ��Bq��y��E��?���!�A�Xk��x��k��y�ë�c��zNf���zӸX&���� z9��[�l�[#ǂ���;�M�W���m�'7<���$ن��1h�ƶ;�ѓ@щ��}a�ݤ�ŕÝő���1�Ox#+��3���~ݨ問8�=A��h2x*����Kh�}�mV��#\'�"��V�w�6���>�'���|+P�q�3�mh��m��zBx��B�P�WIn�r6|}M&(sn.!��Rá���Fb��.�:��|녪hA������1�DU#՗�W��R�ǹvl"N��JD���u�~0	��~+��m��s��_jl�բы��㐃����6�Ru�$q��瘀�^�W4���]GTږI$uV��R���N�h��o6]�����GP�>O3�j�f[T.�|8�X4xk�R���=�x��� 3Z�/-[�T`��M������(I��z�׆�C鱾H:LO��Tr\�-� &� ��&�Z 3S;(}�&���&1EI�(�] V�&$8�,�?kĲȆ�e;c=��XQ�IJ-(^��'F�r���5�|��X3�����'恵qO��ɕ?�z��H��v�b��؞�!}�2�!��y��P^G�� E�bz�]��R2���V��mx�0�0Vp1=���uAQ#`����>8�5��͡&�������Ҧ��J&�.���N6�Ѭ�J��e%��K ��H%DD�Po6�c���b���g8����bl�S��1�	�;v9��+C�~��
7
�`��k_s���oys�A��r�
l��ξ��NK��c�b��\WZ����W��㘍h)��+�@����D����V��u����Wz����ݕ��츣���b��Qz����GS�īܴ��W�T⯉wo��f�%�&I0}��{�GE�+���4K2�R��W���uk���H�.Ug�s�k�(���v�S�]�lNS��j(��tS�v�y�e�ˮ��P}�0�񱆫%��CQD="�Gf5"](mΠ��&:S�E�d�I:���[Y���_=��Z�p���\�k)���.���id���`6�1�F%Q9����bE{� ����H������ �I=q�t��ӄ��'��\.bˀ��L�z��H�
d�zҐ̊9�[������t��՝Z�j�}"�A��}@2�R�z���&l<�\�22��Lzx��]:�m��"k�p;��#<؁�
�����t��V*~��������� d��<c;�\��PA=��	��ex��5#�b�qA����?,^^�+� ��%���)��&D��:��?���7�'�p+�F�i��䛀���?�U���M܀f��.��p4��-���Jdj(
�Wѩ��J��Vh���"2Xr����e8�#OL��0���s���3肍��!m�v�C>�(�	.��P��۬�AJ?��6�pfe_
a�Yۛ6K��p�)�~�C����*���Uq�\ޤ��Ѱ:���Q�2��Uw�Ƭ$���Z��[][��S�8������F��'ÿ�["^Jr�ePE�r��#������ս^%��X -� 5�E�U�c��n����8�
l��^-p��2t t�.�܁�6u$-V	�{�xbe�c��o���ڮO�z*�2��+}ӀiC<@���$$�q���=܌t�K%`Q����-�SC�D�L�f{2fH�c������^t�_�E֗vÝ�L��TY��=��Y�
ԍ��g��vE�z5}nݑ�twUn
\<]lFq�3�}Eu�ra�`)�-�DK�ϔ���Vf��^!:�(��rg�����7���V����wrND��y3u�J3y��dns3 *�}�۬���*�����_N�g'>��7�*Zf,r��m��e7�s{P  2|����s1���#] �e�K�%��:Vg��^�g�)���s
�L��X����)t�%����Ƙ�OH�&<K�9$�'_Y��~h���2��ד��8�?��UeHE:��Oߵ��R^Q�9��8�)H9���-�S��A^�ؔ�@ϕуA�<"�~�}
����r����WmPD�d>]Z���!V����A ̹9������L�5�N���l�d��><�J��	JJ��P�o���/���ͦ��6�}�C� ?�@WT)yئ�c����t�����ǿ�y�!�/�EWr۵r�藡{��9hXI�Sy���^׼>���cG����D�,P�+�
�`Ezᐯ��NF��V"V%`_�$ر�7�Yh���7#�^J�tVs�����W�T�D�6��YP��0�|mO�_��b����a�\��D�
ِ��Z<	^[�v�fL�$�c0�@M]���Z�T���yч�I�6�-�ewlX54zÁ�|�����!�^���
aYnE�*����Z^Pr�XK�@�d�Cj���O��5p�?��ϰ�چ@;FT{��<F��8���IE�υ����C����w�<�j&;8,_�Kr��a���Z�T� ߱P�.�%bҌ7KW/��/�dR�(�_���x)�djӎ̴ݚ.����7W��V��$���r݇� �Иۼf«�~�[Y\ǃ��R��P����ɄzTe�W}�aY;N���zb�ت��/��瞇�t�|�_�V��C�m/�.C�\VB�Q%2���So^΅I���{�;�\r@��%���KT>�靖�m�"D0N��xK�d�݁�a�վ2j���>��w7��p4
���ڜ�ǡA/�gءH[s�tbly��t��|`�O���1i�cbXC#����q��F葌����s�8egʘ��Ej\{m
�.�R�I��m'�<�ow,�!ʆ)����jm�jT�6�_�rr���e�I���X��7Y �e]�]K;ȠC��-e����h��x�����mu̽�7���N��f,���ĄZ���7N? =��jdo�V�G96�uW�(.�ϊ���Zs�p��4�<!�"�<��8��=!�s��A&�/޲�)Iܸ=�sC�H����m���Cy�4T~pVX��6�׳����d��h���mX�����٩��
xL=���j�`)�G-'����'rl������H
��w/m��L�����k��͍7��c�\y�&�AP��z�*b�
'ۜ{���?�Ouv^�f�W�s5Re�~p��B��w[{j�;��z�+"ȋ�ֹ�-@_k~C}��ʳ�Ϻ����8���	ڦ�C �lQ����Ntbc�߲�W&"�l`�:h�"�#��j&�ˊ�T$㧲V6jZ~Ǒ�_b����z���K������x���C���C����⦅X�3)$�z�T*-����X��~�үSOCfR�k�Wݒ����nʳ��M7�w���颕"TY}��!��RZr�>j�n��L�O"����z1����X7�¤ի���a4�+
t*ݧr���M�>����/�*�R�a��C�L�fYj����=�ŵ/���'��Y9�����E���,���9��O7 �4vO�
9V�{N"�f���U��������m��,ĬG�5�y�=��@QW�*n�O��DàX<΍`�2���x���ڒ�ǅ<�P���ԃd����H�,~0�,�!��ɻi9��:acR�:�%v(�QD�'�P��_��&D��h����/����	��ǈ.�s,R��پ)H�jq�W�	H�RzY7_�Q&��#�eg�<�?M��p{,A�Yr��>�g>�yBJ�r�����k��,w`4��l�8��aA���b�B)p8ug��C�v��~C����`A�;�-��w_g(UaD�{��2VF�hX���H��CxE�,{���Ĺ��JU�s>���+.����:�����9�t�W�����g��H����e�#�eC��t�8S�f:Ӡ2UV�wl}��~ѯ���l���B�$�Ъ"���#��LqZs��/Z
�0Z�4�X����犋�v9ܸ���'d2_�wQ�v���vBp7�ԃw�
��k*�o1�j�x3=�0��i1 �Ȫ�N����^2��7�9ނ=��2�$��;�'�v[���{K�$���FM8�(��K�uO�!���{v�Ri_�"|Q�XɆ"eR'(������w��gIAƶS3 ���Wn�h�r$_�w��[�)gՏ�.$'���ǈ��Å�X�39W�>�|���	���m�â��	G#��e��f�X's�<_A����)�6.�ǋ�c��뉠e��s���4��s�$axjM�{n�@�q7��u����wG��	�L&#HNg�:�'����O�2��)�r���5�5AV?�Ά�8Yi�j4���vq�}���=����kN�x}�OuPFl罝�qK
�f��_�W˪$w���Ĭ�H������%'=��>�I?�.��);*�խ�}el䒚WXX|�B�1#J�5<x;��l>�7X����[Q�����RiRU�`Y�c�م.�;JƜ�I��F0��@X!;!�e	u!��e��[�ls�q�| sD�7���n�G\n[b7�TGh7g�vl���~P��O��P��	Q�������4��W,~�״K�����dy�����������KU�69����
��q�����>I,'�B�tD�0>��nM'	�{�����s�9+ro�p�z	^��V#Иv',�/P52H�r�����0敀���)��-�o���"6��7�?+b����g:����F��ݱKq,�G{��.V�8��C�oy��L>��@k��4[@wNI�����7ȶ��V��E���4�ߪ������D�)'���`t-4E?����Ю<;M�Y�:�~��G���sȢjo�� d%��������=A@�{��(ѽp�*`�w�ڠ�*� '�F��ʐ%�� Kk�>p�3�hs��_�_��zgK�u�w��6'_r��5�7OE��0啔���
��=.9�w��V���k��t�w�C![A|�����%^���2.Լ��;g| u��%���ʍ��-� /V�l��e�r(�{�P%w�t�*�ט:E����+�ˣ���&�3��/�w˪�ʜ��O��{�9�b	���c�?L