XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���knX���I�GnIi��Z�
��a}I�~�����S@�*m���p*-!�Tw�P��2���~E=Ӣ��A�V$����~�
�(�K�N��+
7��,��kNg����ȶ0�S������]Ak�uk�6RA\_5��%EB�d 4P���-�,/�2�"i{Q�T��<N_h���k>��4��[0��A��$��Y�X� 5�� �����ef�>J���n�c9�.L�E^�8 K�"��cb���\�V�|R��z+]9�8bj�I�s�w�2ִ��A
 oy�
o�x�>�X��kX<���o�T�Ĳi8�B#aw��F����ɥ^ ����;�p�I��ӌ�I��N)���CA*<ek�Y�r�'��c5u4�̀#�
�3�@�ǉ�4�(�>PX��n�����!�m��XA^����v!��%߃�@tUm��7C!�������q�L�m"R��]Iւ��%#��,X Ami�����P bN����!{�ְ۶Q�`�JxV^_[��ȝ	!ɇ�OV��j_���0�쥃z����6��S�����X&&Wl��~ʭ;Jw?���Xx�`8Y�^�'����p
�{%k���A�>��\���B#N����ߵmw���!φ��OHB��Ⱦ]���@�f~�[*��ف\��
"���躦b�}.+RR�7�����Y��nqA[�'�e�hQ��-7���=�t.��
�$?�My$�ͦ�QX����r�<db�C�a��,��WsE���m.L�~�XlxVHYEB    28ae     b60�5����y�[1��cM��F��r:�N)��>K�ۂʽC�P@x��Q���Z'��4ofbs�zCǳ���|�̫b�UJ���L	��Ow	y�q��冺D��4����ֿU�rG�`�q�;H��^}��z�&$���Q��1���n\���N�����w3@��[0F���sxzIѽl�Aq���
��_*_���v�z]��Ͷ؞��f��UA(�>|P�����t�(io�i�n��Ln�PlC��њ��m�M��7��W/�omUT��r��4.1d��"8�Gk*���
殙� ����5�i�O��A�����f�!$9BA�
�ǐ�F.c��{��T�GPU	Y�B�+�w������][ӻ���D��,"L_��t�4C�LX׵(�j�_O��b⥬��ejOU��������L�tXY��8�D�����DR��۾*�����SN��Z��f��	 ��c�ԋn닐೛5�X�a�<q�LX��Y��U�rao��*Ub`�y��ϒ��� �(HC�� 7���+j�v�KQ�q<���nXsbƬr�N%�4�9\�	�M�C4e���4#Bu	8�Qd.��!jNo�x��+t}j��j�T�էǎa~dÖb�����hjSF�A��( ~��ʼ�O����<3��!fcZl�j#��:P�m&y��O�S��/��wQ�Ťi��-����+D�ү��N�8Ub)��%(K�q#ع�`J.��M)���U�=Y��_�	�/�_�����R�s���p��UF{�ZJ���	v	�.����cQ��7���g%u0��e߫i`��'Ĵ�`!V#n�س�K% ���Cl�იI�ѵ��x�c (��oQb���SA��y|.D ����T�g����^)F�=����̤w��*��*�ʶw��P(HpߏqŠ��O�z��*(^��������J����&F�_8��Ք5t�F�5$��@�����5�a}ь�[�n�_���Lg2�{c��q�?Ͱ��%��`��\Y���Q�C9�!�{�b���2�����t�Ϥ�� ��t��N�z9=�*��~_�����؛�<�������`�#���tR�7�������Vv-������UM��XR�ߔ��Uh�CEmH[�_�hh�ʟ������m��^]ǀ��D���'��[���Kΰ'+o�Qve]��
X|���]��bn6� }��Kg�=�=�dI}��5BȈ���n��;�����:)j���x�d'�v(U��z�3#��-dH�����V|�Y���.��1�cV�%�]=�9 ���sP׎a����1���Ɠ��;�/|��G��y-�����G����j�bԹcݞ��TU�!N .�Q��~׎��6t~�տ�	��/�?ߺ��/ǰ��|G�h
|m���Z��������G4֥-�����Q|��0��'61,{*�&}qwŋ�ˀjh���cO��s������L�ab�J�������)�8��t���C_��"1np��&��L��09�9�;9��3�Ч��
`-�:ɓ�n;J���J�X��o�al'm-�A1��O
�����|Lwime�\� =�v��|�bA4���l}[�#��{q^��a!������Cl�鰼~�|��g�Y@�_G�o�������\�f>Y�)�$v�}�!��*Z�~��#x�y\7��V�)Cؒrw�`J6�^�]4U�8�@)b~�N��odˤ�e��fss#���q�I?�[��RX?~b�W{h$���s�z������n�V����Lu(�3e��?�	� �`����}azZ��6�al��.�4�a{��HT�]��� 5kA�M�ˢ�A}�h�~lA��j�xA)wA�rv)�9����|[�˽�K10tB���6WM��]�ጏ�T4��˰��	Հ�\FfЄ�:c kqH���ݩ݃�[L�3S���~�\��"AE�1,wL8Y�?8G�Z���?:ilɀR�*?P0JƝ��B�ئԹ/as ��t	�EV�dޑ%��9:~H�����ZvKݢ�5��/h�u)��;�N7)����3j☏�<9@]���aL�AQ"����ݔ��K:Ķ��k�.�C&EK�8�'��u�v9͚��î/���v<>l�����EB�!y���=	(��! |3��a����Q����{@��k ��`�	�����L��o�z�b����̬"������5�8���z���#ڴ��:,��tIQ(2�[����xN�~��L�Vp�}W6:$X**֗�P��4���0κX����#��^�s"�{"���)�KR���w"��i8[��-bh(��l�;�*��q���w>"�� r��B�[�ھ�;���l4��] n¯W���5D{�_О��q�B�T?!�h���b�{�$$�ej�b"�`��{4�$�ע�|������dP:��[b	�f�v-���4�|�C�C��i��G����1����8��,�Q�ʽ�����ƒxW���۳����ץ1+!�e�Q��-�~���t}ы�kv�;�+�����Z�S|��F����Z�hA���p%�`�݌�(tQ�lVB��JzZ/~{���+�]����d�F)*���<<�'>�5,ѫ��Т���u����k���ѱI�Wd�����k�1��ck����ʠ�܇y
M�"�̺�^-��j�q&Wp�$�y�xý#��c�J_<�>�s@�q��V.�f�s�5�WO��o[;���?����m���Z���C�����1c�+4[H�Ẽ^�A�Dt�����	N��x艈��V����9�{@�5�u9�#g�![5¦	��^� k�A�H]+S�7���� Z�(�����