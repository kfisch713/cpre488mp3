XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���i.����Sg��>�5&��� �b���7���`�m�3s���:U�ς΃�(~��jEf`��:��4\�^��j�<Cȇ�'cQ�F�	mY���d�q�oq. ɼ"-��@r|I��>�%o[�Me%{V6�#i��5^^�a��\_�J�^���{�D�ΰ�\���	 �R�Q�.?�g�(�MHp��.z���x�uWˉ����$q6�ocbO�sa�d�a�ʊ�i(ݫ`}ؗ�,���+�}(��c�J��I)bB�D#x��{� f ���+EAo��r�������ʤ��M��r�P�6�`d۴ݯtm/�R�S�R�oɡ����s�����Ϛ��C�f�=kЬ�\�=�DR��4ƅ=��dՀ=�
`�|���b(3����Ӭ��n���U�'�QL_'�@o�m�GE6�n^Ϳ��}l�BDF[�TƇ�k�ԩ	��>(`������>�&GV��\����7|uW����t�����f�R��'',-�h(/�Q����M���.{E�M	�r�}�|  n�!��������ǻ뭊/��izu��j�^Ź��.��~'���H�uz9D�����������ԈU�5g�R�Q'�_b�.�:���dH���z�)kd<����
	�\����`Bz[���y7A�gk�qJ�%W��牫?�,��]����ژ��u���Xq�OJIYt,��k"�g�T��"6����j�b�MY7��8���)r�c�ڲM`XlxVHYEB    5e2b    1530N��Bҥ�ON��al����PA�ZR�)�a�Sn5�Z���Fy�L	�K@����e٬�����ey��Qk�\��|� q6F�7A$ӆݢ�ye;�Z�^~ŚWk��,�FΌ�/��U3�����y)�ٕ�ݐ�=��t��d+��L��q򟖖j�#�»:���Δ�;4qo+@r1���6'�UY�R���qJ�IG�.�D�[�VC+'23b�����qKp�4e�7��[�Ƅ}��\wǑ�� E�� u/f?���.���A���e�{�,��6�� I+D������C���	w�F��$�N5T��{�	9��[��PJ��v�������m!����"/7B6�w�>1K[+����� P2�'���9Ȩ�MzNf�o�]4h���6�9|&�-1�ɆO��B��ĕzi|��x�39ٺ�����Hqn��Xp;(a�@�_7�L����|�:x�I�΅���4�@́�J�^���N�_~Ο�]�r�y�I��eP �m��EF��}z���)�v#xiH~h��:V��ǻ�ж�1���bb^����`�:w��.i(��]��s�������d�l�*��V~��U?ط�gZnw��N�r���#b�6�Jh�)>�{��˙x�*��
�o� ��r"Y�]�i.�}�#ґ���c#q$���/=5B���k�2��> 0������߹
��'�cp�����E)Zi�^wb��%�,h��IV�Pݑ���Q�O�f��7���ٓ�[�ʔT+���h|w�ډ(�ٖ���$[�
�q�L4�D��t!�\��Ԕ��Xn��e�����r�nU�Ρ}���w�r�q����u@��36>�pg&�mf���kA�fJ(*���^.�}k��'��y�e[%t�O�늳�|;MӾ^_��l,j	�/g�v���RpVH��0-B"&pܪUGY��DYB�F��	@�10v�vf�C�� �kmh~om��N\��w�B}�"^����N��W�XG��~���/I��cH��|����o�Q���N&
Bu�uVK�ъ�?d�]M�f�{�J2[ۧ��)�T�^�*JQh���d�[�}N@����C��mi��5V���9#ؕ��=����Z{�1��^%��=�έ��d�#b�7�*Ǉ�J�� '�ɣ�9�V�6��#=(�N=�b.�@���$�M"�b�{�&[lUb��".3���̽�R�-���k��A�;�_����c��2��W��V�$0��f��9ܩ�G#d��y���Ą�@���!4҄�R��������OGS̘�)^V�q4�#n���m�F$��p3'd�Wf�!%G2�:`�꒙��(��b9|���u�����zy] �1!��0�ፆp��>�Z8^�BU�2�l���9LGW����� �(	o�q���(���_�a)-�����2п��5mO=��.^�ae��E����3k�Ux�����3���[y��G�n��5u�2>y�n��n
�R��ʴ���0�Z�*[>[�D&W�Rbb<����Ҝj�<��G�g�%��z0�*jeQ٬	�6���Nw�!�XE��:��1.BX���&���x��&#�o�d�Lc�zf�r����P� ����~�􃸰�����9|*�R���#�p�Ҳ�߳ FZ-q�*�ωK�׺��m qԪ�W�����*ٹb�V~Pu�x�ŠȄ*�{K�MK����y��X&HG��O�a�7Yx��ɼ��Ë�k��&�m�l�<�^^�ds� �_"�Y7�L�V�LC�+�Z�@<�w��a�K,��F�]z�׿kW�<7T�㜀x�2��� qIYq�9d���c\\v�:؇�d<\�7̋��LM�o;��|}��(�~	X�1�w��C���<_��S�{�@%}��x��(��R����oG$�$�;��2�ַ2��FY^�d9�y
�i�Bw�$p���-����$�ΰ�S�^..afDy(��]��L*b� ����v�w��]k�GV�8�O=�	�sA��N�Y�}C%���;9���p��$��1j�U��<�L�r�+�G)8I鞣���c>��.P�C{��=����m���^E���}�1	Mn���V ���0%ж]��=C��7��by0Tř�N�L�]0#GHI;^�;@7I�mU�
�e��6�T�S}���^JB��B��u�j��~"�W��c��V<���W�5,��[�:N#x�Y7+�j��p��T	���O�8���.����fC�UO�Za�*�w�q��l �j��!*��
,д28т���5WP��Eq<@'<��hH++�`��`�M����
��B���'��1I�P;�j��(Vb��e�9�9x'����(9��a���A����^h��Q/v��ofɘgn�kq�Rc �9j�a�5U%;�f���#��0t�L6�ߧ���\��~���[�z���p����RWL�q{��}�	VUX��f�A��L"$�Me�����0���.?�kNh�9&������e�c6�"�5�2ZfH�:�ΥV#ÕZ�]�F������FaVT�li?B�E�'�TD�S�<l.��&�[0LXF>я8C�Y��)b�G�&��o���R6 �~���H#��p)ڡ���c�!A��jЖ����������@efqp���$�,��7Z����+/��s��=�0?2���A5�"��>�5}gen0����A�)a@�v� R�J�?��,�7��J-{�U�K�����
|e��8t�O.�S]>��6����v<-��;?0����1:r,M���i�%<	[jL��� ڜ�W���4�K�q����0X�"�fap9���2޹.�m���)s�4�C_���v��*��m�j7J��-;1�p��wX[M�|6�>�m1q�ꝡ���'p�t��	/�W����l�X�S엷,����Ɛ����WG�?��S�����:0P�W�	�^���3�����@�?���q�C�����EiYM��%e8#�)3�"�%+�̳Nm���U��z�Q��2��O%�E�� �',=�R���F}~Y��w�{ʊ;�L���>g��ke�+����\�;fݣ���ع��vn[4��~��ѡ��;�VeJ�&�F�j�:���klQ�	)(J_kg����hP$�LVw��1��I�hA-��$����qF�����'Wt	E�����Q��d=}S,�]<g���Y�3G��ֆ���m@X�%��([�kx`�5b`'O�1rBo���,�-����>ã�~~x�h�&��憘����X��U��)�k����%v%�N���J�T����R1��k�{�_=SXM8ld�?�^���Y,wY^-G�s���t �L�w�t4 �o��������>�����<�����	��b��c�������f(�B7q���J���K4������[-t����?�"�!��0,a�!3�|���ƆG�)�&��ˇ�JM�:�Aׯ��Sb��#@�����kw�!pc[��f�w�y�@f�AX���o���-����ֱ�`���b�H�E����5�m��������JC��C�W�����O}( r9������mLx;�fIɊ����Ws/� �;^�jd%&��1�#Tw��$�R�.cD�~� ��u�Hf�o�LiL�{��&n�rG	��9i�e��I$E��+� �9�>�v�Hn- ��F��y6)4�Z��)���X*F��Z����`�*��C8�e�5Մ^���{+	�mm���B�Y�#����ί O,]݋�����	��v�@��Yv��V\s��	YL��~����a ^�Q�ā�F����t������^��N������L��Mn�6U�/�z�8�9�-�>���OY�p��U��,���f��Y�.r�]P��O{�O���jb±9���~��>��u?���v�4|�&*�ӈ�0"��ٔp�	V=���Ǜv& ���AA�7	A�
5O��ϼ&G��@4�y�����.�BWt^�-q0*F+���s�fx�1��.�Pz��I�����yO�)5u���>���p�H�c�Ri��5���8��ƴv����7o-�Il��5�k~�2Mi�}�d� �Xk��.��KEi힏�x���ǃ�Y�Ԩu��3\�c�����xD�8R�Xb��6�����k�DGSE���҇�X�`������ى(�����Fg�[	�"q�`�^V��g
8@#�����m���ȝ�����wĻ'0E��Dg1N�$*� �p)���yI�u�q��}ц��K^����ǘ!��PC���pW$���(�:_�WN.�r�����տ)��l����I���i�-Ӻ��v�;�䟼h��(�]�?��ҍ�܈]��-,gƈT����&����`i �TC�5H���,�}mE/\Xi#���R��S;wF�����av�!��x��{�� �dA����S��'u!�4��"��������Hb
[�E���Ǟ��M�}D�K?�j:O)�I�aXXE,7���R̆y��c��x���x��Z���~
��,����?�"
��FF!����-z�~q�ʊ����=V�FO.�c#����t�9r��w���R'6Y�#��DƜ#�K��HI;�P���>ݲx����=�U�d�q.� ?Q��Yt����(=�(�m�G���<������"�p��vu�B�'�9K�����u"P���Z�B�����"���T�J��[w�a�#7�ʘ;��E�7(TEM�傪�>�=yj��g �3误S[:�Um�m΍F%뜁��+4����J�|�.�Z�;�A��i��%NҼ\�q�I����[��mx�1DP�K�cؑSav�+iPk�����	��U3+\x�$~K�o��s��}�W���xo}��e܁��$qj�9d��<�mF�i�nDnܢ�*a��1�x��B�OqE?܉o��[�����r�D�Ytm��!k>k��z���P�(d�8)��6�5��d��@[[A���W�$�S���k�A�g�d�j��'�o��V�	�٘���Ac%��e�����/�zM�D�M!���y��
|�Z6�c���6�+�}ZL�D����Zku�T�٬�<(�PRPd����5^�
�oZ�Ѥ�6�=��D6#<~�-�#g��|B�u×�"��R�ǜT���d9>v��s&L��Ǯ7P/9	:�� F�� v��\s��kͷ��Z_�y�&�Ζ-����ǅS�v��uUl��·Ȗ��!O4�?��%�Aܮ"�R��|�v5S�	�-��v