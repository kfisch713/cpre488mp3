XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��30(�*aR�a���W4qz?oF�v[�)��=uEk�9>8��k.��q��R�o��؝�q�DM��%%��c����$�����+�R[�mpT��3�B����/D4.�Q��+T���o�;/
����waå�J�@5[�0��`��M0\�C�����f_X��\�w\<�8ϫ��(�N}(wM�[cxlC�$\W3��ez�%
�P�+:���(x�.ó@}�� ,�}��q�j���d 8���#��j���J+�*+��h;5$���'FG;�KueΪ2/��9�O:�ҋt�ػ�f������f4bQ6�7���>�0}�&���,�?i�%fk���5�'f�����|��	b" �A׌�_�0�a G��*I�s?�Q�h�͓���d������%��;�u@ڂ�s�8Fiʿ���z�4 tCe���Q�F;~�P���[��ZkӾ�*�J~�V�s��5�͓��sF4¥Y~B�C��hݵ֙�y�$w 6�M�����%��ˮ� k#�-� d�<]K�T�ԵQz)��Վ�R{�G�СBր;���{ 4��_�Z�F�xԵ��
Km���a�Y:���d���Ҕɥ����]U:˚�: �)�[��^�=��3O�����+���QH�3F�O"�(6jH�PϢ}��qE�>��4�)d�f�UTtDHɕ���q�8�T��ź�{6ۈ���E��i���bi��j:n��5-���qm�� E	uWUڛВ�3��R��JP���OXlxVHYEB    2326     980���RM�?���>'�'}���7н�9��ԕa������}j���͔��Dɔ��Ӱ~6�Y�b��%sa'6N]SAkб�MO'��Fn�os�q6%��U} .C�k��v�7�Vͫ���A����B)(qU(J)�$UZ>��S�%��H�̅X�����p���V�ެ���4`0&���N�z�6����m�c�fI����9*+G>0WnY��=�6q��C�3)l��!�,x�a����5r��!��xի�g����Z3D	�F5��@v��[엗��'��r����$QVک�rAi�@X�7�hC/��6%�d�v��,��Fx��SQ%�r������ ��]��6{ٖpe�,�����9 0�6��毜����
�Ί���� ��ˁC�r�uOur��1By���`��m^ 7i��z�����u�L�+��ea@�~�ޅr����6~J��c��,���+0V�|-�t�y�c<����g�\�?4�\a4踬���I��@�"DKн�s#jͧ��u\j�e�N�w9\}��x�������4��ʂ�ߎ��Q�g�M��x��T�R����.�lc�!�t��{�&��X�����Ն:��,�}��q\;��,nv��6wǟ��l����9���$Y�&R0�#��B��۲͟��&�m�K�rO؟tɼwC�d����ű�v>*�uq�&�� 2���-��o�4J���z[��`ޚ�m�L]�0���S=$ uowl�OwD�o��+��)��2Eo�j����V�q�L��BT�EUm����u/����d8���- ��L �R�.����B�vi��Y�H<y:��]�#r�Yy���#3L��>��'���km����R�dK���:lV�u2��f /Z��y�@H�\�]�]�7�z�Y���T����E9���r���|*k�^�¥������/q�8�����\�g��C��W��C�����RW��d&�4Μ���ȍE�}�*p���ȓN��QY[v����RM�vۥ��Hj��e��H�G2hz�����l�k����C&:ǩ�i���\�߲q�,�E��� [���)��d�e��QhǮ�'r"�ۏ(�Z���Г	���G sX�T���5w��p��u�\zvJ��aF�P����ׅ��b"?��4�X+��G�{�$����E��c�D�7�^�������30٠�(�"��k4��D�?u��4iRr�w\U^=e�K��a����0sǄ����{�|^��gfo�:�a�Ƞ+�#�Aү�c!6<���MtOD�&����?S�R�= P������繳�62U�H�`̵O�`{�T���L_���EM��Y��*�+��dՓ�)>B�n�=a�}��&���1WB��Q8LhWTb�L�Ǖ>�!��S^��^�Z9$��
��Uϸ�i��I;FS:Ś���m(�j��.����8��Qf4���-jJa�GZrRk$Kk�2i��j�W�D�q��{Ƶ!
��}O2������X�L]������
a *r��\���cF[�zL���=D��2>��7p�CH�$v��5Y�n�K�Li���1+��Lux�חC�g�~�zk��T�˅�1s ������^�VC���m��ѧ{.oD����N�w�Z����[���Fy�K��4Vޅ;0ۮ�����~��� n��id奖�2s"9B����*4?���tb�����e�UB��+�R'���TtG�F������V�Bߊ��Su�5ܳ�`#{��߯d���=&SV����N0�GY<
�r�jӮg���/K��Y�������s{�<P�t�j��-��>S�'��,�~��UФH�n�|O�W������m��\b������6�N+�M '倊n�\��aÁ��RU>YӒ�(&塎%3�o"�F�J[���0wAH'�3nXd#'\�&�#�2����ݺuy��ݸ3
�G��������L��%�����Q$�L/���7L���SΔ�H���L�>n�e.v�k`9�Y���� �s����~��j~,�����	GF�,mD����@�}�j$��75@��H�dr������l�d�ԸG�T����p|��ŋ��]�櫜R����ߜ\����/�Y�$��]Z�4���(v�ҿM�[ȳho�1:L�GaO^�ś|������Xz���S�]�iZ��:�]�{`�N��vu�M�$pі�����O�j�m����&?�N0k��B1��$5p��*�����T�^z}_��wF�tHGT݋�P��B{w��A>��y�(e	;�]���w�����	��R�A<:~���.�� �����D���z�V2��d�L��