XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���1=H9� Z���~Ħ馦����..\��d�l��_7/wa7����.�+�߲}q�u�t}j�C���b��&C VP��M%G��A,�D/(ز�W�B�����^�Z�ԡ��<ѵh����щ5n����D��q?�R�.P�� Ц,cD����d��e�г�Bx��A���ѫ����Mu������;|��wS1���L2���>0rhwH�N�{��9�ҽX��[ 1ڢ�4L0�szZP��{%~��jytOW��Y<��!�[� ���;p5�U�y��GNl��ڄr�m�t��!?��,�e���]�BD&����ϳ�&��v�+�2�)fPAC�p�3�:TN�C��+b�ХG-��69�Ϫ���]�0�R+'���f�г�D�%�t� r�ª�ؚrBp�5��맇c%�2�ޞ��yE� �fCe�̵�fm`�u���bG���rU��m�jm�;)�r�22Ɓ+{Go�+ gj�np|�Nj���%c��&���j���z�6JR�_V?��Uo��6���w���,���s�X�Ac����Zfo�,b�&N�=Yta|�F��f1�={z«n�٤�uw����-����-�J��:_;#蹞��:�ËBB��M���㯢���X^�`§+��9kv2r�.�.i�����(2�O��\wt:^3d� ��~�t�7!?��ܠ�Y�����!逍�_��퓳��b4��|�<[/��mY�
ҁp�VX�}nXlxVHYEB    15bf     890���v΀h��;��M��QE4"1��Ms]j�1��O�T����,���iY7��ߠo�(��L��,H�<?��h�a
 �%x�Q˨���<b����WT�zL���|i��a�@��tD��%o.���*��}*�rc�����?K���H�q�kW�난()G�odC٪��<���&�/4�Ct��h	�È����L�Z��R����j[\daP^b�s޵�֞�B�A_�:�,���Ҹ�����S�0E`N��Eֽ&��a�5��� 9vh;��LEm�a�&a|<�����[e>7�s���;�ȕ�m˛�H)B�|��FZ)�A�r���]��:֟��e�Ak>�[H/�֊,����@�ط��y�Ǥ�XzNG�|�[E�7����3�۞G̠V��%��J~-�qy��-,�ş�G�C�劧?D�C��tG2]~k���qk�TD�j#2xTvI�3�U�}Ht�9�6��!�L�o��� h����<�[��Y�"Y�[�ܟzk�p��t�uA�m�0%�A]������I_`��m�n��f�����
,�(��0UD�	c*�y�}x�f����ɖ��tv#�%Hm�<�`��0��k��][�HE2�&{W��G)��J1kӎ�.��C���GX�eO���#Θwh���{wn>�ҔWK.L%�K���,l�.��e��ߨ�) �A�a����y�*ɊQ/��k�R�Ɯ�6]�����g�[���xsU��<DdKݍ!	M� Ձ_O*	hy�ܮ���[ ��	��/��"�w���ۭ�Єf%}	rR�}ZX�1p�(S�AZ!���;�.|�,dl�����7�4h��W���8�"U��Lsfu���`�_c����w�����$�L� ��|��{ې����u�a�P䚺F��v:��%O:em5����Pbt�Fʚ?i��ȇ=����|.��c�~M|
~�r����jaD�TJ�ݝ��8f�84�\M��ٰ�bM�����ڕe0�Y�\�:#�jE�q�y����D������wL
���q
����tS?�M�l�~�W�6��s�Н�R�.��˛d�B�\���G�]@/־�b�{J2H����G�~U�MR��N�&��1Q��Lń����|v��������, Kk.�6����uԡ��uT��_��~�H�X²�-�r"I�Wy��\�v��
�\��Z��{�j+�k,�dO����]�%�i�6)%����d@���S��R~3����� ~q���ŭĚ~�Z�{��J���`�k������W��@������wh�e�[
�˂���Ч���k%J���N8@V3�����z�#a�X�LnJp�	Q�hK9��X��� x�KL�J��CX�d����kh`1Gz�v�U�ތ�y!��R�{=Yt�k��z�VG��GS�i��yV0Йy�Γ]v�?�g$��|r�k�倹Vm�\� �O7�V���2�_�R��[࿘���dQW��`"\ 	K�n�B{�?'7�ۡ��.tޙr�w��~	lUߖrI����ӥ�֊H5�D���������[A�{5��@�J8��:�B�\��R2ұaW���}=��2�6�ꈢ�(�7��se�9�
 �f��3M�Up��&:��l�:{����o�l���<���Ix�yʔWϭ8�'��l���g�q�A�n��v�/i�s�/��^�?O�p`c�����BE~?_'��3*х�
���[�a��L��<l[�����s)��J�6>r�&dK�:�g���Z��yi�Ow�|���2�"
��&�~f�����*P�|�8��s��q�@7�QĒ�n���N�	�d�dQع"B9�R1��Х��3��QeĒ���P���29%�,��l�r�I��*��NH�{0���������J5�\C�)O�^7@(�o��I�@P�o!t����?���9Ծ�*����Y+�4���v�%H&�����J�����j�s���|-V`4���(0�I����q�����+DZP����+� n{&|������T NR���~BM��|:?��K�	��<���b@O��bQ�>�#�7S�H"ߙ��$F`�셺�