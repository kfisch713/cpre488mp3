XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����.�"@��E�tQ1Xm �O�ZC3�v�M��T0�J�26&��Q_�B�7/bF�"�9F���<����$����U�&�H�j	��_ ]<&�Q��%���L���T٘}}Rx��ٜ5�\/n�o��G��G�Ƴ��?�Xl0�s�	}�����z�Z%)/���TʬB���͗����;���(���S�PM�ϟ&�eX�Iʟj��j[٭R�ys-s�3�ف>�ktW��-/��E:E2&�5a��N@��W42��Q�9E�})^M. �"~QK_�*��8C+��/bs��Q�̖��h��(Q�aI�E��K�Q��i5b� �A�U�k��܃���`��,�*Y���b ;�2q�l%�9 L�f�R���<���Č�:�>��{��Li%�3���Z�9y6A����NV�ʔ����w�N��29��n������d�'[b��Ǯ�~�<����]��=�$Q�׷����l���(��
o�-�Q�7�]?}U�=p!��^���6�����(H��E��1AwՄ���qL�.M�Sh��<1u��'_���(ݩ�Tٴ�]-����0�7ܥ	:d I}��IM�KH����o���\�G��	t2.��`b��I�3�^(��t����q6.G���GNB4���1�M7;s��f�E������?X�!�+�cz��Ɖ8�ŷ+�!�\�ZX�-G�;�H;Af�T��.�!BI�j����&Me2N�$0��e���Θ� ��XlxVHYEB    290e     af0e8
��'�e��L�n��˰��m�ح���C:�1+��u��?C/f)��*ts�vZ�"R��tٺ�à�ڄ����M�Y م�o:�ىm ���>�\5�����$8`�I/[e�G��z���_t{I��M��ʢ���56ܿ%�lO3��Jg݊�T�W�C�Zyg�L
��g�]L#ꓣ���/��Csj�%��!�ӝ�h��X'	�U@�yހ&�.��y �7�!���3���e����II����d�0W�?:F51��N���Wr�k��1@�,\�p��U�4�k�FW+ob��sc\|D�@���Ȣ��;�2��)k G"^�*�uW��KK�,����m�M
jeCV���+���>������CU�,���hƓ�֩�kެm�ӭ2�%�^{���q��9������8=��$��2�%�luSѦ����5�&'�-������)�}�K�-ҢQ��@N��+K��ŗ�A���:w9[�clʑR�oP�q��U���X�,���t/u��� �v�Vg�Y�4�lW"O��x��}��d��Zd�I��o%���t'�)NAFcX}�E����>M�i!L�]�R��y��5��t3�,�y�Y ־�ͼ��A��Տc̱�ި8�Ր������K�]��=P?m_�y?i\�T0a	��X����t�� HM"3i�4�s���^2cw�n����Y�5��u�U��\4��4���gY.�d&���-� D��`��ǉ?��,q)+B~6g�\a��:��x/uB�� ��@�&p���̷��>����C67o8��U+^ ��-�"u�,4zpc]OɃ����ONH�=����7yaQ��+S���<[�->/��|��E�?~�b="-�DRE�+6��.>,�8�	�7����V��}K���^	�10a�(b�B���x(��A� |��ZO�|�����1J=V��n����	���̼�WDmB�E����/��5�FR���3�:����9@ൿ��[�S��I�w��_��y�0:~����OD�PB�u�A&��謒$�VB�wӯ~��5��{���B�|�AD����4s�j�+/�EK�J�J���w^��9��ݸaW�c]�g\J,z&�N84K��Ȕ�@�2]�S��?v�.�o0�ig�I��������7E@r�,�p��V�c ���� ���vW��9�I%~��"��3��G--�O����H\�e~������K���ϭ�X0��~4uǌ~,�Kֲ��pe׷L�;� k����|�Ef��\me��Y�/=[-:��z��^Yƙ��_�=�b\�@P��P����U��}��
��4F���<k�<c��1���D��(��j��7�ِ��V_R��Bw�#7�1F�J:A��?SĈ 81��'�#.4p���J3�P@ܽ��Bg2"�BZ������C����
��!�k_�k3�.&�U���d�SϚ�:8��LOs�0J�a"��S���O3K}��?�
ԡզ�\Ǧ황�+���Ǜ8P�9�����c�E����r_��{5�~\�O�+f�:�Pw���&�-D��j�v[��ƦM�C�@��U�:I��Ǜ�";�?d��K����Sl��&|�$B;��&D����`^?4�	{5�8�W�9 b=X_^>���v�u4eO��H^�g�C��Ulb���1��PL��5̢A܋�Q��0���1F��j;ۘ�#��4�?c��~�*j�ؿ���0ٌ.���F��25�z1��(�J&�ԣN��,% U��P0���z�7�'�Ü������������<�eX� ��.&�tP^�f��K"�D����v����i�S��8y.�Ϳ)���\(p���,5k�\���,X�M��c�C^�?�����%�ox-fF�;�dT� z����Tb0�!���'�9z�`��g͂�<�[���Rh����W�M�^فeS�NH"_0���]~�S�e�ƕ�������Z8c
�0F \GlN�p,yռ7��[^��I�����8y�؍�8�����7w�r���"al���s�-�V8��_�u��i!"����G�Q�~H\���n�`$�q8F�o�U[��`jf;`��
�`���m��D~7$�\ą@���Ű������6�(L��Z\y�m\UHL�T�z =�1��U��jφ|��[[�j��$e�'�\	X����.ֽ���]�~��#9A�����߅/}ٖ������C(2#�-GO_�U7ysm��?ZlO~&9q���QfFYuE9] ����b�c����qM�t��D6!���������
(����x1�4g�ݗ"��{�8h��t�~3&�zh��+�[�?���фF*�mv�U�+��1�X�M�;�TH��|�p^�3EqYE�G{�����7��]}�آ���%"�ƛ�;�KF��6�U�����	��-Aa)]�2�4���t2Q��]�S >q@��p�V	��P�6?.\TF��ub��@��R�����o;|�&J��j!����09sF+PO�zWjt�����2��'>�̔ql�X��j= �/�e��#//ز}n���w���8ʋqȿA�M��V!L[���X/�������vȋ>~��7d�����u!8%Z�J��&�$S�m	1r��)ZD��Eܘ�U������ɦƇ��Zc��Ng�h.J��K��ls-Y�9>_K�3��n��P�Yb�����rť&����M|P�?�!�b�&�