XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����d�>��^�rv�*ќB�ּ�A��U6k�03s;L�<��v�Vx�p��``�
��h��J�q��|���=�����~��BI�����f�s&%C�&�� =�	α(�ܿ��ZҼ!,L�,(ϑ��O��1gH���6�Kj�E�+��ivdG��5��]�o5���<�U�͚�q[�E�<o>76F��QT��4����rFyuS/ģ��gC^\�|��X�it���ȱ/O��*��i�6d:Y���0�u#]�\01�΢��<Re������E��L<�<=z ګl������A"�4!��ڹ��s�d��N����Jb�H�&;�� 7/���5z q�[��2�Nt�y��;�Jɛ
ٝn�^�>�t���^䊛��y�܀��[
���Z;�^�v0--��۹�j�oi�M�C�;�,�Vil�D��ǝ�N9!2��{r}>��[wK�)MwzVl�Zp���#~r"B 	,��@�N/�{x��Zh-��G��(�q\��ya�2�,�%�5�l����ǋəo��b�=��Ep���}�wB9{��v3�Fx�;	G�~�D�t'�-���tڱ���ow(�3�1�2�X�{�|̂^�{��s�V�����@on����m}��]�B1�#� ���u�l�XhH����XS�,u}|<��n���i��7�T}o��zS\�������e���Q����;�D����������N>��*דtm(�J��3�?��$;��ʶ�VhK�1M�XlxVHYEB    2b39     b10��/��ͨ7Wiȿ������c$�O*�Bt^��s�����Π҄f��[ъ��h�Qc0Kj�\���iv����(wS"!�	��艽�+�CrGj��WΆ)#���³
B�����R�^��ZS��S�^r�������6��B1I���5pr���q�/lW������l����k~��6���B�S�D�tn������Q���q+���iT�yv�3�b(_�̷8h���wg�`��\<[�)6:���t�_�GRhZ�G!ߧ#Q���UM=
�9�F:ר�����
�cJ?,3�.��*�񸤪~C��x�L���?������{<-�X���tc�;�R��Qa<�VkؘJ]xƠ������n٥k��B�a���=�LͲU��<��e=ZK+��C/�%�����StC�(r`��1�L����5%�ҫv���d��6��|HO*�R1�#U]qvS|��X�Ʋ�n��YѺ�����ˮ}��y�_�)M�.~��>���Q�����kڴg���-���.i��q��^)����D���z5��Fl�H^Ɠ`]�  �[{�1���	���Oo!��5�F>c�Vk92�����h� ���U�~߿�P�:!�6�Cկ7徔ĺ�y�F$ �C����:���� "ϧ=�`2���[��d��6Vl��������t�9�J�"�\]��A��T0� c &P�3Xߛ��9�-)B`�z���YPz4�.s��i�ԋ�u-�����~�m�إ�G/?�X�|o�,��<�7�n�0y�����(��Kk������E��Z�3dQ���KV��oZE�e�<����8�J�����]�U*;�q��JWJ0a	�N�V��Ӂpc�ɯ�DU���M�:fGx>�5�����>H.��v9�>�T��T'�گ�6oB�]�ϭ��2���yA&@/F;(�G���!F���r����Ph&�N�ȒΕ�ӄ�XO�E��'R|u����~�� |�Pn��$Ef�`�?�ʵ��IU�L,��p��-��T�����V�p�����n�)y����לfW�w�;<|g8xN����:z!Ο{t�yp/_���C���r<�Qf�̹,H`G%�8�!���&�]j*��Zpt�5��uC_#LƜ��f��6*)ޅ.�����"�|elO�3��V�OT߀P���L���Y��F)@����j�<yD���#=PT9T"�^�%�n���z��E��{�u!1��A���#�4A��#M���},H���;��y�Ӽ�{}�$۸z�bS�=��0�'.�
���Ɠ�+����-��؟���*�Q}l�7���]�Qr����n�̧�E��F�^ۭi�w�N��,�ڒ�Y�-�x�Cd�����s�\<oB2�'x`\�{�,�Jy`���[n`����:������	:V�%��W�Ϟ��ܥ��	q��(fsy��
;5v#<�����:��*#�%�:�����3�4���r����%z�G&��5��Ww1�R�Asc��Z��O���H���8���t�s/5L����%��8�)���a���!�JRN�5��?U��P,&�g$��k'p�,{����t#.�,��7\ܵ�yS��[���|\,��㨗�*\�+�1�x�s(k�!��יj�(�ט�m�P�-�oձ��v���o���C硐~���"�t��5�$A�{^�U��5c]>�RL� c����c��_Kޙ����L�ߞND��y�C�a��Y�'�1f@H�`�oZJ�%Ze��� ��Y3��)3�o8Cǻ��Z�+����ϡ�| �I�����ªH�δ��E��"F�( �h���~M�V�!is����A�5X��	i�v�)����%��$2`�7w��		R���S	a �t�W��-p�_��6�/���ܾ��.���FK������;/��!љgX��69�V#ƣ�b8�Қf�b��k�׿Y���!�eg�s�Y�ҝdzP��S�=>��������<�u�Υ�t .lR����	E#$��Ƶ�S]��%:� L��kb*�ۯ�ߥ�sD9�č1i��P��V�<߲�2�asO9�^$��B��@��x���?p��1����ٸ��Wf�ECy��y����`�7t��Wd�4� ��$�8�ɲQy�E.똓��W���3c�CF6�+ps�|�R3(�]5����ل���
�`^ԩ��/5/j
[�q� �Y�SQ�5�|pi;1אN�N���1���^t���v��G����hwՓ��o�Wea�Y��V-�<@��R�4�������ZS�DR���۵T�}��MAG�t�m�荫HiO�2��"FL�9Ca��=�N�5]^��ijȁ�n`��M��Q��V�0(|T�DЉ�-�5+���vPFv��0���e�nǬS[�M���1z%�J�0h �G�����W�_>�w������J���f� beB�k���7�Lh6�&P�,��ʔ,�a��0ʯ�ڄ;r��
��lN0��-R ]�L�|�@�]ؔ؉�b�m�]��. ��d`�0 ��dk��X!�!�>�U���@��I���x�f���\6Dü�9��׺�zD�mg�>�f7/--��k��E�<�B�M��!zۛ��K���:Hl<~*�x]I 7��f	��~�ޱ �$���%��4�g{6���߬�ϓ�a
��݉��n�M�^����������ơZ����Pp�h�H������.��F�_�x)�M���c�v�s8R_��{#G��&�W)��)�+Bv�騶�~���Y����0d����O���a�i