XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��xM� �p�I@���_wfyn>�I��J��v�W�����l�,���<����L�Q��^�[.�$��F��8G�"�һ�5�Ixk��z�����tc#��k��Z�����_Y��[�cb� % ��}�g[���Q�h;*,�n�$�'��6I��#*���[Q�������@3�e��CF�m���>��]�Fᥩ糧�Vr��]�����ߒ�u�M� [6���%�$cE5��	��.����\"����v��kT٘�����g)�&N��	H'{P�U�V�#_,�UrU"q�#۳���[�3r��r�$���E�Gc^�d!t�4���XMC�9�I�2$�:P�B�2�ؾ�
��8�9�>-=N���F���頒я!��M���N��#�'����K5�E�+�B,�J�0�@�m>��S)] ��'f��L/��J�x�a�@f C��#��_Kc��c3%�
G׊�y����̋F����|�HMа����`GD��Xy��,��݆�[L>E|�����������^ٍ�ܭ�O�}2�/�#!��'q�4.��D�Ѵ�'`CE מ�$��6�ɷ�qhʇ<�Z�]�ɺO�c!�=j��9���J�d���-v����#\��x��p������f9�#S���\=��	���[.��F��tE�|��98*v��@�y���4����Y�m� O�}5���R�Y*��s��:����3V�A*���]��-P�"?+��%?t�j���8ǁ|�Jڵ`�BXlxVHYEB    39de    1170�����c��}�gM�]/����	��5�U�v���p����~{�:��7� �耡�]d$�LP�:c�v$!t��B�ws�:���V�"�����fLb���#�a��5)�����̵���]tkE��6(B���j��.��:���_�
A]��o��
Ým8sX~���tw]�ߣ�QXȀ&G�6�������h��q� �E��g^�Ւ½�[�֏	M�"���� ��\���Yqh�y�:�͸d��ۃ�0r-��O��w�l��3�x�Ɏ�@KR����6q���j�H���48X�m�F
�;��:4�~,Ԅ=.u����
�X���l Kx4�7;�/B.wk,m�ߛ4� �ޝO0��hh`˕�A�7{�*�������C��׎��.�����|�헪��gh9A��9fk��!D��ޑ���S��x����{Y���\7s�48��0���Aw����?f�x}�܆a:�1���T��%��Y+�^m-� ���-��]�~Q�
FfŚ0���E��:��k�X���І�%w [�������{=�Z��[ ܠXW}o�&X�KN5Y���K����ȅ�ֱF�.��<���S/�Ѯ�h���"��z
�wi8[ѵDI�G�6�R�P�a���޶�Y����8ψ����R��*�?C�fG�9�._ ��@�����Dp�!�}C�D�%��X>3f�V���n].y9����@	�&�4o�i�@��E�{l�ߌ�y�TIz�����m!S?e�s�"��s�ìfI�m}��qȻj��Ec�0s���IO?�I�qž�:�4�۲�>�5G�B^k��D��-ΒڔG�s���2}ɟ6�D\�d�3�f:U��u?B�����Ib)7���Lo4�c�#,(/�Zka�g��sm|w�Ձ�|��i!�0s��6���(Gv�ѩ�e�BN��쒅{ǭ�QSC"��2�j��0o�/[����xN��8�M� l?��ϒ�+጗�����sGb�f����՞3zX�y6=>�G�=��'>f�Q,��g�j���Vd7�,�33��K��J��ɟ��*��|�i�Ԕ����j�&l,L�HV����Y�G�4�$k�ݿ��)�9l�	����`-I6��vns������C�b8�yA���b��eFo�:ߣ�� ?�@�4�0��!X��ax�z�S:ə�)>z��#��R�3��B�Ïd��,��
�G���O�;l�^�w��K�=�:C�|7�7���[�AO�ꝩO*���;r��I���X�I ��:さ0|U؂�Kj5��ƞ�q 3�PQ(x��F<����Ju
�E�g��ʗ�ٖ!�
H$5ټ�7�D�Y#쑅��ގ�<%�X�n��E޴�V��c��#��`9��U���"���4/���}Q_^"�Ӭ������[�kQ�~�e���������J5 ��.���y��dG����P̈B¥�3R�wFU���ebZ���jY_��.	����W1�|����Fq9ʶ�T�D�F�(�e
$���W�v)p���Ӧ���?�΢d����՜�&	���(뗆��'�o�S?g��9��p8Yç�܅�O�T-/鵪۷)��Tw��u�w��}χ&J-��|x��%i8&�ư������R������y�Չ$
�Sy�A?8Hd�y�UN�wa�xJ�PЌ���bc�0��1�����1�<�C]^�X]�E��
�M�_�.g܇��'��&w\z|AP������}�x~y��6��V;�I��6{ܐVY,��'`鸑bͬ�.A�&�"ryojF�"C��SP}�]Vf�O�9pw4�Eci5}�A�����y�B_���S-QsJ��@+�]Ñkv�6ABI�yߜ�n]p@�uPQxA+��o~�J���1^� \-�hb
%
2��7ru�M�,{B`���Z�R��+״�������	�,S�z�u�Pi-"0#E77�l2k�ME1��0��^r^�i��lX^��{tE2�R@��WqO��/f�������Y)Fȝ!��OHa;��7�r�0���)}u@�x������[��w��=	@�K!�p�͏2`�gcs1�4�B��#V��h�_��R\�{�`��3�	j�����&�?=�R�������v�h�|綴�0dz��B��T���\��� '���tڬ��q�h��\J������>t�x��b-�7b�b��6�|�0��T"+��ymtT�V%(�?8O?tT��m����N���U�
ԇ=Z� "!���d�x�Ae7&<o��� 
A#��L�DM{I����4�8%~�v���Ń��|!7�Ҝ�ҩ�YAc�9�m�Uśa�	zt�%[�=�+��Z]��s��_�i�}�Ka%�Y\�#��]�As�H��~�|��ΰ�����Uqe��ƪ��R%dQ�Ikz�׬�d���R� 	��A��3 N$��rͫ�p��d!֘SY�(�1�����PY:�/�;�o�6�/#!DmFt���K6-!H�'��M�E���45��^&J�s-�i�Y�R��Q!�Ze�F#���4C�	��r(g��s�|���Fc��T\S�����u�۾��L_�U4�E�`�4�V>��1�(��5E[�T���MIUG&�A���(ꩱG�,�O��?ߓ�^��aCM���ӓ�-6�Y��]`GVU��li�g��H�Rz�F�������>�/g�?���T��Ǐ1���;m���Kю2��	kw��=���-��TI��ľ~���ͣ]F��xHvs;g�"�1��|e����Osm�#���d:����VxK3�ٔ%ԙ���aH�Vn��c�.��x�.��`GS2J������&Q ���G `��Z�0��w��>�[���h� :�%
��H�~%Y$��h����`E!t��(�S�� �9%{��
��'Q8�6��-E�>I���s�:�Q�qON��31L��ܭ$c�t����=�^u�=�k^�w>/�Y���[R�Ő�F;��=s	�az9�*�+�z�5��o�L޾i�=_�먋�OZ�-Yxaϖ�B���E{�If�z���ʡ9*���Y$c��2���_�h�Pfy�En�R�b�sY;|@\�j�9H{�S�-O�r�.��>'��# Q�%i�K��?-{����]Ϸ伯n�fQ=Yz�FQsϬ�L�t��!apOx�Tc�GUm���=L�]5k]��S��ZA�R�����5�l�U����eoK2Px�[ $=ݡ��#�϶��靊qEir-jX�Y��O���_.����c��;��C��[���l[qk��� ��C���um)��t���wF>Q��h:�h2T^��hvt�'d�vS�րD����ۭCK���F��'�3yB�m^6� ����"s�&�T�N�с�+��T�P���Dx�m�� <ތVy!�u�z{˖�,�̞'d��[M7���&�������o�O�A�k�+6�Ŕ.Nk��M���b���(� G�ln���,��a?���\߄�߯;��2��2��{�="�r�!R���Fvl?�A��D�J��O�������O]#뾲r�R��������! )�?��*,�,�Y�f�t�ɺ�q�*��}�%�"Ί�͛wf�e�K��������C˒3�#�;�iS9]�HS��Ts�����}v �w~����p0k��!�VA��H���Ȣ���
�E�M`�J�:`��|aU�g����ja�#DP&���������#b|K�a�3h�x��z�휖0�F;&H�!��	���Ҋ#o��-2-z��cuHe;:��X�)��q�E�� %�zMEo�x��`�]X#Я
�H�0�L �tݐv�����*�?G�߬���"~��ɥ�+?�jF
���'�-�c'r�4�9�ܷ�G��K�NJb��2�|>��W�6�����2�ż��td�.3~D1�e��xă��2���Nǜ�;ڞ��lN�h��$��>����fe�OI�)�y��-l�B���Րf�4b���3�� uFIΪ�Ҭ�
����%��7>ٽ��k���U���[���ZX{	�冋���;y�Q9H*�x��dт)���n.N�h����<�*�g.�o6�u�!�L�n�^:�N�/�v߱��W�D�{���@dE��7@pһ���/u��잩���fs�=/݈�I�E{�P�WG$P<�������L�TٺC2��Q��J0.���2�䉳��	ͧ����ڦR�^I4q�UD�����x����НV�2|/B�X/b �voӘ�A�b3��c������lU�����/G<Ѓf^zOwmKH%&vW�!=
B�5����%�u{��Ĵ����gB=����1�R�+���d���L�[�ˢ��#�*9?�u>�: