XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���]�����$T��0��}�a�ݐ����\�xT���}���SI�6?R��b2�cq��}RaT+K��ؗ B]s:o|�.�k��tK>�.���h����D��cG��g-UJ*���y)b��'���/S;����H�������ZwX���^��H�m�;v���_7pS����BG#���$�*F�U
v+,�5�'^�61,5��:���I,-l��h��$�=s�F��e�5�p��5v`­����DJ���naT�{VӕJ���Lf��߈hh��V�I�t''��rQ=����
Sy�B�W���{�[.  �1iE����TK�oaj�KlA%X�=����Z�3�̩f��e�6�$3���e���Ό� ��7��.^ĳ������%#v��H��{p�Wr��Ċ����#@� �h��K �?� �J�����H�Y�����^aT���'Pd�H:`�K �Iw�2v�?U�H8�刕I��H���پ��bܥ��<��绦��wθ�=� ���)r�'O�3%HQ�`�)��m��T(�%�G������I� �G�ϒT�6�٢r֧���J����v,�Z�P���6��|?��x\���	5n�%Qh�����?h�.��֮�2��M���~
�Y@R1�'�FF�sF��M�c�������E�T�KR��8�T�F�6�ݑ�<A�������Ī Ds�^SS���r`ں����,}0�o�F��ȸ.a%��-
��J>���Z�k5�#L^ئ�XlxVHYEB    5224    1740(� ҢK}A�k.?�a����O�E
��� �֗O$(�?�УL�E'�G�XK�5��v�4�V:'��]�Vb�:��eq �I;�Kkr+���A�Bp��<�b*i"���hi͛�}�8����"#�=h(l�\J�A�aS>��uS�A�<��Kz<V��fW��s����r�$!��Z��/O
�y����u�"1A
�m�r�� ��j�n�R��*�_i�.�s����^是OMbA��'AM��;k�8uӡ.?�Y媗>zx�1��S��r	�b�4�+%
VѬYCɱՎ�e_W�y�W�6	�c��Hݻ������	\p@���u�C]Q%eR�b���>-Nz��X����Tt,[��1��bieD�V�*�&�S��ZJ~D���}����S�$CW�����h~Ν�j�_��{.�;6k�z/�$%�� �7R��_k4fg|�a�X�$*e�A�|����7�PZ�ۯ��X����e��Ł�~q�(2� ~ݽ�����M��ςހT[9f�b�Wg��9���#�đd�� Y�}��B��"F�~,I��"iNW°�Re��t��B�V`�y@�ӡ=K�/D�Z;�� �U��Ć�(c>��h��3����>�O��R|'�탎��6^�]��Mߣ� ��*/������2�A�Y績ͱ_��k�W���º����hr�^���}қ�C,�����e�Uc�x;IiI�X��r��y�y�9"D@�9�������v[�T�\_č���;9���@�`w�`<�!L�9J̆�}� �UH�54}����^��gē�\L̖Ѻ<��x��ԏ3�싖{*m+v�@4��"��^�T�c%!��g%�R]�:(u�������T�𿵏D� ����1m# ��Eº���C�,β<ғ�f�
�o�+sv���b�^Y̡٬vl̰c��O�m��_>K����~�9�?-�Zn$K��VU��kp������� 7R۾�-��Jt'l�x����Y��H���-K�r˚`�dN۫���UE25;�"�ƚ��=�%i,�>�F�%!^�&�/L�����B£r��V�Җ�?����,�2I����ꢝ��~m�p�R�x��%�0�w�(%�C�hry��$ ��Xў�-2��r��e�~�,4����+�����n��4<q�IH�>�V���p��Y��O�ׇ����J��zψ�"al+V���v3^�3�C��e����6scmm�=�w�\��oB�����l��������AV���h�����h�q�2-2S���5F��9�T�|�K�=ﭵ��$������X��8���s� 2Ζp��Q�>S��*��j�ܔ�I����K[k�<��x�0�����T���!���6�{ϋ^8G������fHou�> ��<����͉N;���Q����|m,2��T:���<���]W��n5�����\7�p>�U|��4e�����F*���po��2�+YF|��YG��^�2wx���J�M!Q�3�Eyƀ/rO^hx�ϜߓׅuB����[q��6ȯo.D����v�h`H�2ؔ���ąZ0�n �P@��"%p3)�J�q��й����58<������#j�  ���rۮ����!*����=;��P��)td^��q�C|�	MU=�e�g24X��pm<ۏ"k�!�l�"	��P=��_�KB&g�S`�%{N���KxN�(��>".1�x��3P��ϋ�m�Ģx,+<��:��q��b�f��(#���8��^���?5f���Rp�n;�� ����������U�C��9�����G����~�*�̋�X�s���6��8iT���ef#y�����X�����U����`�oR����PTxH^�{.]�PG�iA��	ȼ7aP�$��� ��oꌗ�� �!�̚A�,��$� ��+٩��0]��Z���f�Ô�TR��$�(#�̻�*�oЦ~�j�C�f����B���m�fd)��7��y7�p���ׂ�3���a�)��%����Z��� 4Sy"�4Q��j�9G���\��˘6l�9_o�S���2�Q$mw�� ��B�n�	DN?//!��T.�|�1F9���n99*��{�*�i}���u�&�	!�%D�9$Y�dN�{�t1�S���c�,�I�Yq�D�8�V^Y�yx���0AɔP��! �3G�\��As漼��E�ٝ�1�Է��"���t͂�����B��%�A���[*6x��A�łV�s�iW�9����Y�2�h8����%�ʘ�?��<�b<MPr@_jg�MvhX��WH2 K��󐝭A�C�|m����z�z���ph��2XC�w���Ո
O�|�@p��f���1���K�ws(@it�ݭ_�2�1%�6�3��2�,K���8Q�a}�	���!;I�����O�F@2S��	����T�υX9�}�+�Oћ)O����y�NB��q������{O���,H|���Z��f7�ES?O�$�;���P�b�������V����]&�=���S���G��1U�*�c��F�f�����`���0Cgx���l�h�*�6:���-��3@��x��1�x½B�m�j��� �1Dv��/:b��BAb��R����Y8'OF)��f���F��r��`�'u�	�(�9����g�Wp1�\R Gᴩ��GC78n��5_�3���|�&j�g�����,��R�VP�{U[��7��Z�X�2vomIQ�&\-���C��������E,g�+��w>��g���n����x���;p�ZG�jWu�W�V����C�*$c�/bL�*��@P��2ǜ._��o��6�kB�ǚ��h�@&YN��.�^�W�[�U���sׇ��up>9ЃSx��e	;���q^8C#��M�D��* ��].{�ō��]�
��>;&U�ճ��91C���9�UB��~���� ��H���M����XuM�.����7b�ղ6�B���&�Q��W�2u��=������.c=��1sêrM[��!5��U��!�t8�˕�ԧ���m��<Ə��r�� >���T����y��f�ua��n�\	/
���V���-�� �6Ak9�O08:�K7��h��M���'��
h!��=�	ʩ^
/g����^ذ$~g������+�>Dơ#��<�{~�� VY�����j��ڎ_��S�|Z#�[�`�\[5���W f�E�q�XC�����SΛZ�E�N_�_��K×�.Q����eρ�|]�ʬ�L`�X��� ���S�O��t�T���5G���a)r��{ܔv�vI�YK�y����;�d���5�[ٌ$�Q�e%M 1��:�B�HC����*�
1�����I�#P~:����ڪj���p��X��u��j4�R*=�
3�Nf`�l|�% *�.:�W��\B��2 +�m2*�s�xU'hcܔLj��abI�Q�J>�_=���1�ݧ�O8��D�3�������mʿ��<b�������XRO�.�ãF%w4 T%��kVY�9�C|I�s�����dj��ӠJ1�j�a]@��=�2����z�Y�X(n���R�d5��o7c�}Ec���Y��K���~��Fj�s��UB���2���e�@����T�xJ\?��t�HF�����nСgRE|ì:��-,��C�d{8�����N��j� ��00b�A+���k˺�h���� ek��[�>�K��n�y��E�4��0�Ep'�x{ſ=��>���X��z
`��>���=��{F|�b��
W)��S%��nq���G�稱��UR|�q���պZ��[���RE��sQ�}:qY^���u���]��0�šG�1�=��C֗�U�j��{�l��H&��U��l�dL ���p?��h<B�g�ph/�<��*#���e0[~�ܺ����\9�)k��ԧhEn+�^�W�Oû�yN�-y��~��Td:�� ��b�N��
����@@�6Q����k���'v��wf� ��S�K?�\�z���$�t�q�3�2�_��
�djo��u��'�^�y�+�� :b���&�j[̿���]*�8X4��	˕n���ShQ���]�r��0��cC$��>=�)�Ė�5.��"����y�Ւ���E�~�R_��z來x{OAg�N�J3��踓�l3�V�1Yf���6Z��;�m��jǷ�<����&`*�h���>�����
����g�sbn�'Vt7�[ON;��p}��w�&����D[B N��U����n	���UT0Sp>�ylP��g�S<�T���$����=��p)����γ� �
Ì�c�C~�N����;�c�����t�� ө�ณ轳���dk;7.�T3�F���D�4��kN��Z����ً~��9�q; n6�BI����N$��.�CT������Qw`�H�.(
�:�Q%�)�����&Y\~h���kY-s��]��h-9IC���O!G�2x�*Om(��?y����;-AU���Ȟ���3�P�n�.���l0��mkY� OB�S�g�yH����j� )���!��^��ߑ�|(d�\+X1��hX4b�����9���hn<�	}�	s#w��U�:��j/}� tZ?��a�2�	}>i���|��#�$��Y�w�� ��5��Sn9���EZ�X��KK��f�ci�� � O!�"��/IW�/ź�~E�{�����c=��(F�����*b=؀���3/>K1?� ��&;����M>��}ʆq{O������sh��&���]p.�\R^�|��7`����g]{J�L�,���E5-�����4`_	ؕ�s�W������~��4�X��4�+�!����`�i���PxcY��eϪ�t"����)EA�h��8�q앿��S���P�V���΅d��sQ�"�m�X|�X(S�^�'ܶ&{�g�v4���������ѴFc�2$�S����o�k>.���@� 2�PF�_.P��� �tz܁�<��;R������(��Z�[��iW͂�8=��uh�":���z��Qu�s;�+P/�	#�~��8��q�HîJ^�
BjR�� �k��T��Ø�i�}lC0p�p{���SD�^�32 �t�	o��Wc�)�*ut������~�L6@2�.v��o�Ǻ�;0�˫��j���<ơ?i��[�8��:6.ے���'��������?x4��S�l��P�dA�o�Nܛ��:�Є�^�rg�e�#�n��M���g�1?�u�}��)�'/y��ޝ2Wh��{�Q��S�����/��%��~�X"��ɭ�Ο;dM��aB:�s����ӂ�5�h�G�њ]��]� ����o��`���nU���\��3W��L�Rm��3�9�y �-��x�X�R�s�om� ����
?��b�:1V�eS>{��D˿=e�`9o�H��VcsAڜ$i���u��~o&N������B�?�w�8R���2���;�j�[�bZ\d=��޼)r����~��]h�����R�c�bG��=��7b>,�<c��"�ʾ�G�x>(�~%�f_vu5
�ԉ�^a����3z������yj>����G6��ϩv��j����O͙�^v"҃��r���P���k뾤A��(��گ�3�쩵Ւ��{��e�\;��"����ͭhmEW��ݴ^"�\�#Lk���
�R�㢿��JEי����t��y\��N�UQ�D����� �D�g�m�`sV����ê�'�*�4��u}�v�� 