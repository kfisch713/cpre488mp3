XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��D���F��푀���ܮ����#��:K_��5[�4�!�w�]\���iF�q��R��)��	3 �,_�A�@ijg2�bKD�>_J�7����t����ކF�~&ьID,�9L>�A�7<������@�S�Q��9��r;mM0���޹-wt�������X�,��'�!��Bb����c�Z�V�6��e���j@��_n]&�W�C�\�A�Dr�ul?�%��,�#��|4h˴�)H�IG�Ǿ�.��
���A�c�nJ�W���߫��bϖCVf��N��#
D�o�v�b�LB+���[ѓ�8��/��)~������߿W�|�`B��? :�a��jsHYD�nwB��Q�j�8�6�v�%�{=��E
$��Aܵ��M���Q�����1�[�J�",�QJF%B�.�C�x�E�C4�l�l�$��>`Sg�������.̞���ͷj@�{ol0%x�W$�𥠽�x��:i�3X���úB�,����m�"?�&�c>�u��
�56Bx5Q��o,Л���V�V@��E]�@����p6���Η�r��s/!p6bQE�*��,���Dκ�w�@��%���,�/J$Z�G�v��̚�!�Y'7'�^��t�9d��e�<��m��V2����Nx�ŋ���A���
Apx��` �򍷄wˣ�䏗Z�ͳ�à��}�4��Ii�&t�'�M�-��U�G�ųbQ�0qip��`
�u��io-s��;�p��q���nkP:�WD���@t�CXlxVHYEB    4052    10f0x���$���6��S;�P���L�m~3�|G����C�$ʀ�<T9h{�Cg�5E���V���������{Xb�qA<���Й�i��.�dԗ����B���s}dN���j��;���1������p;>���ڌS�G�M�㝗�9�W!d�P�A�x�ۄ�"b9;8���d���9����>�y�i\fx��"'Ib�`e��,T���5Ss�� 73�Ct�<� Vv���դ��6>&���|���z_I�^�h�'�H�7�p��D�̰�?�%��i!r���˶dZ,���Td�rR�I�g�QYv56�1R<9�������ɗ�9���5����L�s���Ń�sᓣD1&e5�޴�,i�ɛ��Y����KC2�:E��V�����Wl�Q�]�l�Nm���ɖ��6������grH �v)��t��hI�%[�՘wMe~�-��#a����*r��N�q<��䳆p�8�� ��t�ջ�^%7�Ե�6$�ǄC-2�eAֺ�R����l�C����_ڦ��t��rz;$v8�ƙL�&@�ɖ�;<�u\��9�D��"o�z�| h�E�ks����̀�#�pv��
�yi���T������m���-���Ԡ�j~q��(�kJ5����6�s8`,c\J]6�����;�_p�	��8��򒳨F�գ(��v����K��Q}N��:���[�E/�_h�����l�x���P�e����FR��Os;a@?�o߬s�ڬ�IN�0�b�Ɵ^�6a��V[��|���M�����C����f,j�V�&��8�[Sn�ı�dW�#J\p���8��q�4����
�Ǆ��n�e�D�E����s�xA�M9�i��'��8�F ��B���):Y�u�� b��t׾}������GC˽��u�� P��9�`����S����01Đ�����W�y�Oy�t�1 N��%�e� �Io�4��&�&_�i�q�c�
"��W¿Ky���[��|�wW�ނ�K<��S__L��Q$H�wM��%d��i���Ց��v�xp,^���L�R�\�$9zzT�GTM�Z��n1>����Q��\t�s9��L0�-�ѕ��3��(�R�9��N�EM���HT�a��ؖ8S+�5�'7`���>?�S�rf����{f:���펫��F���5�qs�Kq����b�ʃCg#�1J2�`�3*�)�c�|�]?�XT��L�K���s�����p@i<����� �ħ*'�u���܄v|OqJ�����#a����Ѓ���F����D2o�k���pa)d�
)�\�E����٢�`u��`�p~>��#_���gZ,m�O��ل�馨�4�P;��P}6�U���*����أ�?� ��jL�P#����J��F0��>�K�r(�1|����2�HH��F�֮ �T��J��Qͤ"l���S���~�SIZ��b+ՙ�g
8��Dg�p��8
T���9��,�[�O��J�}�Oܽ��;�x�Na#�S7�����,f'|�.��f�l��W�E�eX�n�@��/��Jv��!<7����u���)||���E`X�ϭ+K^�2d�ҕ���A�C�c���w��}�]�o/;����$õ�B������Kh}> �/�vJ��eTɀ��з��B�l9	!|#,�f����U���o�ip��P����vF�H:lE��몀��ܠ��*d�C!�*��ҭR�"@Z �=�Dd-��6�z��|a�ƴ
����x���p'�]��s?�n�Fx0!�+TS�:�1%�EmΘj�WV�Iꃮ��h��7'��}!��\�����@y,4��n`jm^O؀p��V�=7F�6ݘ@E��u��՛��a�#����l�Thq�'�<RF�"���MY�	����uK�����)qZ�rҼ|ev�e��D�/�SC��<qMI_4�[��7EoؤQU	������Õ3&ˌ�~83g�>�zK�e��U�9^���ҕ,�V:�)�o���2r���"�Pz3�Y�����W�/o���Z�T�����.lX��-~t$�ok^9�Y����
J2S*g@N��%�9��v1�km���Zr�' ��N�W�E��+���\� _m����:qA,H��m��F�ʽNL�ox��'��.��2�+�~��Yx8�z@���C�������(Q���n�s�K���F����tr����5v�D @�����OQm���D]�0J'r��Y0M��� ېn�ŐXcA�O���h�Ɍ�g_"}��{��+~Bx63c}�i�-8�&B��������C�/o �k�$<R
��m-�a~ȑ)�1 ���5hX*�f������s"�
#(:\��yq��t��N������J y��9�_ۑκ��	���i�)�U|�x��X%����j��H+Ov)ey�B�<�=��X�����_���w�p*Io�f����<�9�ޭۗ� Jd�-�	�W��6�d�o�� ��tUD�с�}��0F��]������/r-��]��8:W"o~zH�|�����x�<�l8�6�S�12J�X7����wVgg�`�Jk+
i:�߬�����~���	@�f�)� ��U��O�q,:��e�  ���>�}����}�mL�O��Mؽ����%��>8�7cM{Y.9�Z�{7BX)���}=�Bzh8۰�+�+�Y:�:_�P�M������UI���E02������v8�ݽut�s��~}�;�r�['	�������ۂ�����Q�W���$��-j�FO{�y�n�~��D��?�B��un2�������@�>f/`��4�\�z(�	5/Pe������ص�,)%�O�d�gP�s���m︐���plj��x=n��)��_a�L�:�;Z'x�F$W�q�A�^M�Zp���J{�ns����Pg�p���s����.��;������8HN�|~�&�S�֦;����#���nqV���H���Vr�ȅ�sޠ+͗ A���G=8����J�W^�J�o��y�GQ�@��#gIP,�8�8J}@OJ�Y���%{��PQq]�k�
衩�(t� �%_�� d$-���OfNC���y���!�vӗo��DNX��_s�[�G:u]� t>v�A�7�k�Q��*�f���N�i+�+˘��
�_8V�~�9��%�S�i
��O��k7�ֵ쩫P3Z��S����fx �1��ge��1�ҽ�|�b>]�l��h,��d���Y�}��IEM|��WL����G3�C���LR�w��s%�h�܈�7�jAƥ�J�w����6�:��tm�6�A:y;��-��9
T{�/?+o����d������g
��B��.��FbRƝ.����?�:De�-f��M�����ÊŁ4u~�������̱�M*C�}!��.���X�� ���+�!���׫���6����lf�gۂ�g2���ky	F�ǂ؉F��U�E�,<�_�tm���v3a��r!�6�m�ҕH����6k�ꋁH7�%�X�?G�T-�]%�T�S�tam�(�46��WZ�ū>ާ�r��3�zU�&gӰ��ƕőa��x�9��z�r���3�Yo���W5k=��Q�Rd6�ѡ���Y��N6�|�@�K?S:M�'u�F�\T�����n�9f���d�;�H_� �T�j��It������]���B"�4y��krBG8br|�^כ�c�+<��Ê��/�'`��_g����ԹV���0�4���Ɋ	5��,p�n:�����JЍ��s<�dΚ!�I_�����z�6|�yq�T������?������q24�xnd�T^4�m~R�����{gv���Ĩ�,(�B�w��Ѫ5�k�^��u�t��q�F�?�q\�
N<A��=�I��t'U���yhV�z��`z�7:>ׅS�!2ҝ�v4[�΢Z���j&	#W�O�j�xr��}�v�Rx����j~���Jt"��g�w�h-�4���Ekq����t�X�q�e���K�⣘*�x��F�3B����07�N�aS��kL�#�K�8�z��P����]CC�E�U�t�43$��sU��A@+7��.W���O_Ip�4�բg���:ڳRQ�R,۰\c3�F��|' Su.劈ӯ������"q����Ll�`�\GT��	�	k�SE0��D=6�~��4��