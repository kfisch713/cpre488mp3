XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��_%>��Ik�'l���{���sJ�O���/�������?�Xc��S�٦C
���D���>8�
J�Dw�l�%���(Q�R��l�J4����4�Q%�A='`8������4Y������S�(�kQ�'�0�%�&�L��q5��G>ʀ;z������-s"Ȯ9�*�N^p�[,.���cU�o���ʓAE��[ܡ���D�z)��1�`��'՜ч�4��A��3פ��hщ}��cch�9�f���b��b�6�N:�W�Pd��!y���3�[����p6�+yeG9"N��و�n*���4�ڎZW)4G�21�/8Ѣ�ޕq�R���9@�������n�� D�L-��z����NNw��d:m��'��j,��q[:8�\Lɋ���?n�p��
�cg������Le?CVg�ӊ��#7r��{/ ��3O�[5A��j�C��\�?9<�틧`��J��4M���ZR:���1�<b��҆���Gz�ZIa" ����r:J�s�U�*�w�u�;�4��#�@qU�S�~i����k5��}q��v��)����ޟ�8�$���23�>�)�
������ݾ�Zz���D�6�_����|�Ƃ4���9�Y����_2�V����՜퀞�^��DZ˛�k����?z�%��;e�hQw��o!Q%opB^�4h}m���(�BQ��s�o�kg�nA�LCx���V��];���>*�<h�K�ׅ݈�?#���ygXlxVHYEB    13ba     770���ZF�pR?��{�$��}��[}E���D��u�F���p��&At�c*Zp^ڌx@��AF�=���Oc��U[��$Bac3Fd�1�ʢ@<=����0j�>	�趆	�����d���>><�M,� %S��9L���X]���9[8B��U�v����6���j���m�kȜpˬ�'d�9�&��!Wz��Љ�e]����l��Eqʧ(<%�Y0��z�����v�c���}a�]�z�.�Z�\�\�9��PT��F�9����0M(h��7*����\���D��m�̭���[�9H8�#���Bo�����D؎�56z�%� ������qO��Q�)���Z'6/@-�u����+Op
mNx*:��y5Iv�Gn�m�~�?ؤ,��{��RPV$,�^����6<2����>( ��.�vF���vM�~���L׆i�@��f�����J>�K�P]�\܏�E!hi�Gm�n�����?�xpA	N���g�䘓?}O��΅o�t���l�F������A��ع6I��;Sۍ��&;c72Z�M��ag��{�Ic;~k4�������� 
�X����]�'%P�su��+
�p{VE>A`�j�!�%ŐHSǧp�ޣ@,�t}�I�,'�|��Y?c��2^U��|0i[f�|(k�����b��	TQj0���T�y��`��<�a� �	>���|��8t|};5�`�ǿ��+[p��9�!�<�h�����S��X����_/��]���eܮI�iuZr���?�.�y�OO+����%�=��0�r�K�Q����Ր�����hF5\�SS-��GB�m�����x_�Leye������͝�`���fu]9S�@ԗB?Œ�61$T%�V�?�R�ʿ�[��:��K���UED
�ϸbπD��ڼ��6N� 4��;�����+��@��

b�%��`jy�&pAm�g�^�Jբ��dP�&r��l���9&+��8�mM�Y�e�0�~V�i���b�E4�?� #�|%b�%4�s�*$rڎ��-�,������։~Y�0��d��R��^=ք��]����#�*�
��Ɗ�T����i|�a�t�Y��{VE����&
;į����Ƥr�y�g|#��>T�a�+Q��Vݕz)�,Fo1|I[u�f8&$y���E�n��ND:���`���\@V��v���s䊩�@�����%�D������r���8��m�l��7�<��m4ߩ�B���G0����˛(ϕ�~�ݑ�2�'�����8*��Y*�$zm�S�C������P�	)�D�e�4��I�R��'LV�U��j$լ��p��!u����?�,�{��[_H��n�m�R��&c�9O���ڭ�T��Y
��t�a-���5�q��W}zD�od0YD��9��0�'`�8�3����3�@�oU=��#E�g�gq����.|��ބsG�}�;� ����k� wq�w'�{����
�DD~��"����WM�.�E�|�nφ��\�<ʶ�1�cJ*/��p��x-0΅��gh���A�����V���G��l,��c	H;����h�I�Z�����Lq�Y�aE��(Z���Zl�)��jm�0���n~X� �'A��8�	�z�6Ej�4'<��Z=�Ҭh�V�	촽#�#;��ݵM/����`�/A`CG���-5>/7K0Ve��T��?������Kj/��5��ڴT�0E��>���k�ۿ	�f�
'2��;Y�Rf\ZS�fƔ���m�1�>'�"\�I�U��ڨi4}��O�b�ӆ-�I�N�P�9�4!	��0`:��m[��~��>[/Y�	�1�=���4�#����ʉ��