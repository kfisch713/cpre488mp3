XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��X*��2z��g�� �8�$�;��#\�Z�]�~���z����V0>I�-�	�1h��pfrl��(p��G�/��.?��;�m�W�^s�s�)����.k�Z��¸��6A?@�A*��@�3?s5�@��l�m¥�
͕�/�C�j��\'s �_pݛm��i���"[@�3q��F�ܨ�o"�T�Q������B-KCHnz�ƺ*�;�u?�
�+i�g��%��6lF�Zil���J�@�j��c�����R�=fH�/vo����:�&Ľ�
����﫴
�]�I;��O��U3(���[���
St?�z�)��3�<-n����:4�4������ i�	��û~<��
j�i�b�߮	U�ƙ#��4`/J a�	o�$Z��5�5�9d΢D/���aH�P)e3���~nP�x�`Be.�C��M;���X[3_®�_z����'�`�J/���I|����T1���G]#��4DvA�N|;���(t��z��Q�yF��{P8���S�4��<���3Q����} ��0\���'
&���W` �|L*� ��e����_&��͸DDH���efk�a6T4d1qIj��g�6ʨ?tMJjFy����NQv���O�^�]��9]+r�0�(T��݊ a��W�����YA�\���A�������C�aY2�($��FBv��o��MĐ<"�������F�|��^��ٲ�[k��(��My�?s�[��[�(PR�F�IcO3���!.8XlxVHYEB    893b    1e30�����a�CgV�g��q��f���@cc@���^��%�n�oB���ؑ�w{������l�U�e.�wG�~n<����?����3,'Z�Ӂ�W�̷��;y/~��� ���L����	��ȭ����wh��0L_^���I�b����
��o�O��1�;�	���α�)�������²>,"�&;�N�tG:L�h9���I�N��F��D\�� (@��P�P���j9 ����lg��p{�8������iJR���3^�������t7�o�������5��{�%v��^3N�=:4Q�{XR�Xt�w�a��Lj͆��@Q�OH�H�F�<ZĤ��6���z�ŭ�S�$�(Z�mh���Q�c=�B$`�	� ����}���)�~X�L;[���t�E��
L3��s��b���Oms��RÌ�C����>jB|>&�WT5����l����%��`�'��S.ʧ}�w/~Bn��)�V��⼅�g��P~�څi �³HdN�dZ/��?O��[[Y �RBz�:�a9mJ�!c��R���,����9\§����5)GR�R�1B�w�T!]t�_��T_�6��.dP��f���U�j��
��7�����b�
u#�K��۶K����V����&�癞�ɢ}XF��.�G���㊆I��Om����@�G�����}b�8"Es.���	�D5~_�lk�����m��ϣe�NOCPH�w��<�����-��g A��qѭ�p��mc�Vy�F����>��6w��;Nr��L�}�+	��1KEK�h���#|��ڍ��T%|��/�Ё4�Y-J{�<�*r�To���E)����'�є����2,OMB��91>4�Ǡ���w�{��vܟK�Zv�~��T�R�%�w�'+�
�2�c~迚1�BT
ǌLC�R}sx�K��ǩŨZ�z� {�vB���4%�V��u��W+T��s���Y��U@�H�Gk٨�[s���r:�?i��i�Bt�IV�t��ċ{����ȱ�a���k�Z6�"��q�Se��z؈�5�C/��5� 0[FA�b�m�C�3�N�s��� O�ضA4�n?�r�@g��M�����O��߽�i[��yt���!C�7M��HKl��f0yA�p~�F����l��aK3@�wk�+@[<�&��YmV�j⮢��d�Z�=G�#���|+}�*ݾt�+r�C��2HP�S�y�*���(��ѵ���?W��:� ���H8<���U�{#�/��He�#h�fF7��0X�L�?�C���3Z6F��+�п|�!�Y����RS��r�'�.����A�)?�6k��y�"xK|vG��l���r�M�"zo�OK��q�0r����s׵�Ч���^��T]C=3F~}٪��)Y�F�>�5_E�b�a���+/�(�*Z�Ic>,Ls�qj"P=:dԒ�"����$��(��G�[C6�B��.H��󱅢�[��Ƕn��JY�]���?�������&��^��ސ�$�F�_o�"�>�ٽ�u,h>���z�n�)2|&�@���3'><��.��~gΘ�t��P��7�۱��u��PCF,qy����&�����������If��5���:#"eM�����e%��dؓ��;dg���ߪ;E�8H��� ��z�-R��"�ߚ��C�u����"�l��' O^�l�Ej�����$���>��.XϪ{�T��"�k��B&b�[��w�u?�sIђ�/���g�y�}�'�7���i$&y"�Q/�G$��a w�O�Q��+�@�'��������Zf�y�r�B�@�N�����@}��hVM�I�5�p�d�C)����GU�������Hz�ΩM��f���5Ƶ��n�]�g�x���6�x�h�T�H>f��!x.g�^Kŧ�"� ��)a��6��������=K
�lt��Ej�\����:- a�[�@�n�E���o�%����%?�H���{�B��˼*�At�|��|���|m����wi��B[jx�>/����?�e�������x�0�G�Ø���.�gZ[����:-�:>�#q���� �8�	����[�ǯ��U�\Y.O��� �}i��҆xr�P0��Z?=��~���"v��!��R죬��Q������P-�-T�����l6M9��F�R���ѸZ�%H<.�]L9I��:`��Cj� SLZ	�n%���i��6v�������u[�ȻHD�t�K�`�8���?iS����Ġ'T��T�]D�miA���b}{S����b�X�'a���2�اix���9`y��qw�x*�?����8@��4]��Q�N"Pj��[�ם8��rM���D�=��w�� �T���9U+/-&�֖\�GL�^V�\�J(�g�5s�1v���Xi�=-�w��T!��"L �7<{~�����.��1iHLۧৼIvn9��PnT�"��^��K~Z�Êc\�B,�C����=���>.],�{�]�c����tNx���E��`��
.�o 5@��(s���[����	(�.�t�T��K�w9�So
�Vx o|/D$�ƪ�~=>�M}!�v[��(}>4Z+���G+�:b&����/�Py���xb;V�=˼�vh�8,X{���f����f���KC"�-�#t���D��=�_�%�|H������<jE�F����'&�7�d8KI� ��P�����%\����@E����B�UtB��-���MU�}�	��N�LcT�g�l�����s��Vl��f�#	����� X��t�n�}��=5l�	E���#@�AN-U��5��XV�t�x�-�F�+����}ĚA~��K��r�9�`[�6��O�V��|nHmΉ�n%c�-�y �I�5$Vy,ԗr�ϣ�5>�[S�)#�>����w���]���"��'��O���9��Ļ�"^�ٻ��$E�wQߩ�y�W}q)�n��}'#�&1Q0�p�q��0� ��?�u�Gs�7���i��<��P	���������_ʱ�,���䉇!9'���v��U�l�|����)4'IM�['���� {.�5��/� �&t���vF�_�ة԰rpUU.a0�f�T3��(��_N�7���Ksh*�3`�xY�y�e�20�1��ӢR���vć!fQ7�؁M�I�G@���}�T�!P��qڦO#Z��),�Ä�����Fݔ����O�_�x�^���#8���	�&<W�o����������Z�A�Ln�$ꫤ��Ǿ�)E�٢C)b�'Nw��|ˊ~�D�b����겼���"��o)���z�;&M�~���坱�#��a�k��}#�X	��Ѓ�]A\�ɳ�ol��~�p�v�5)��s��K'�S��hR���"�±��h���2c�걥/ �}?�+�t��b�S�d0���M�$�j�>W�;��)p�+�gGl��m��̠b e2��zJ������F
6^�DQ����@��Ipq�>�9�V�qm������q,�P�,C_�Q,�&6l��l�k���(��nb�����u�oE�~NJR���we�m�C�vjQ�x�]{�MHFѴ�< �9�n�z �_�����V���-=N�n��!�N9����I+|��NOكw������1}���'弬�>Rᡌ�n��k�E5;��t	c��1�v��R��:m`[3��>��Zt..�|&����ID�`*?��ƆWz���8�s:�����]�}���f�^�5�lr1×�'nYDv��Sn��/��CRc2"�a8�� ����y�f��#�Ȏ��(v�tYg����8�A;=̣y�"�q�Kt��M7D��%�ռ{����S9��F���#��@3��E_�\X��{�M�n���OdN�5@Z�2��P���^�@sw��©!�KH~~h�Ԫ�3k����'�HO�.s��f�߼S?����R?����ޭ�*m2"2|��$�md`�c��a�r��<o�rt���ؽ�`�i����}?ѬH�Jb�7M��g?KyH�^C���&>;R��B��j�y�Ȯ�"�u�Ak�,%�u�3�)����2�`��}\�~SGEG&6��7�Y'�
W&��"��a*>���^9�SJ)br���R���~�8�ս���t�Ա��&EQa}K�K�sG��\��dSPI���r���
Ԙ����E
����:3�a~*��0�m_dɧL��g�ӊOd�Y�F Ӿ.Z'�y�L�"V�*|�5�[�f��O�(#`����Ѡu۪�Iq����.�hн�v-	��8I��K.�+��/�]�U.3r��4�� Vd�k U�u��U�ի���'�x!�!��
�+�H?��$�&?zwr�I�Gn���/ĥ��D�7�c�F�>N�$UbA��-��-2���p��{��O������L��Bݞ㭖��R㾪n�Q%37O�&���JP�39y��sM��K�՚";�5Մ��G�l!9�X+L��C���͒�U(ֽ��R�n\<7 �F@���T��̰�!���n�r���Ӌ��xET�����ΓD	���2ï p�6� ��[ԏ[�<Mĝ gdT��fj��6�s���z`�o��\�Nh,�v�\m�H�300�,L��TVdT;/���#�4Ew�0�c�3�|��s}�QY���i9\��oL�����(ibw��+W����\�nq���!���Wܝ2��ݽ�З��IM�N���h��MB�'!#h.�kp���:��Ӟ*����	�$[���h���;T,��!�-kH�ao�Q�\6�z���9[0��'`ѥ��\�;-SV�z�ElId}�"��b]�斪�(��eA�D�[�.L��J$�X�X��tݢmV�o+��MGHX��-�F�<.���h���o�^�:�D?k1oo��2D�r�	���2 N���3�AZjb���H1�4cR��r紿��a�A_�վ����6e�q��
� �L��[D@V�g���R0L�*B�Q���V�rF{��f�ڞ�69�r�C�D�J*XA�t�����({'W����O�n�nzj��e��#$h����?�^��.:Z�>�.9Wd�k�3��h�Al@U�!���`	=�Tv&�A?a����q�F�E9KS��ߟ^�2�Wgb����C�3�fw����EŜ8�T�|?`�c�����;Ȳ�gT�J�6��`=��A�+��3��s_���������C�#��à��{gZ	��uZ���/�(�+�����	�Q\!@���'#��?[�*2P��T3��y�����y��o�Pd{�w��[���mq+9P���NrB3�i7KY��'�_g�d�ι��޹�8���(	�̜vx����d�����8a����,�] a9��9�Br������Z���FA2r��u�� ����閛�L�{Je�j����\͔S��#�4� A��} ���̿���NtӨ�8D9��jxL��v$K�zrS�>
,¶���6`�7)x�x��%�t�aId�)�{}���IP�(~���df)_��0=	�oN�F�!_�}�Ŵ|��-+�*؟��c����\>z������o>*̗���x7~�Jj���r�����W�{�m�}���~�M��Z�N6��]�S����te���{O�Zn<�֊�q�Aؑ�<�	2�����N���2���O�����u�-
&��*x��c<nI~�Q8�&�$C��1��f�I�1s��0�
�����J�AB�Q��` ?����=>��"�4hz��[H4���dÔ!.���-{&�7���S�%{ԃI�|"}E.��l����=rǬV�#׋N����ȫ�w&d^�	��'���P��_ٍy�W�Rڝ�%�n�ks���z�Hˋ�\{��$T#
�SN���}y{"f����u���a���=��u�{wn�g�|t'���` 9��R��ǩ�I�91��I̽���)�Lk���Wrl�*�=�
��Tm�q�%%��[-�&-e����Q-�%�5\���X���]h�kC��N�F���9α�0��W��=��TA|��('����@�h��%M��Ϟ���b��T�AW	���WgT��l �0fN�����[�&}�:�˃2��p,�a��aTr����^��W���̯.�"Z�r���[�^v��V& <�S���P���G��rD���c[���像�9<w}��qW}�ow�w��z��J���\z�ӑ�F4���y�?I�'0I\���e�3V_01]R�^Դ]rs���_���Z� �ʈ��[ƉR&���j����^�ٛ���g���Y��{��PW�h{�T\�# ���3��'5�*\|�p�&m�]��õ�I���:_DF<��S�IT���8qD4��,W�y�m��|���LPUGR�4�#�>�[IE��},5�E<�U�������4|�D���2rc^.jOFa�t|�]N<I�pY�߱������(���e,�WAHi+�P���iw������]n���@"/�OLb�y�J�� ��+5Q���%`Ȳ�iK{��Y�i0܃3�^��
�������.��Ɇ�j₤����r�=� ǹ@�����W�daW�8Oymw���[����h[,�W�x��Z��rj����b�����;s��]A�\�����Z��zH���+���y��"��FV�}�'�n官CQ��N������ogp���μ^��_��g����K�����q|��x��볅��tua�)#d�^	�P�u����j��i���hN�~�{�c���ӆO�����=�ޓ�rR=��]�M������M�����MZ����"H�Q^�l����������c޽7�����ҭ&��rC�\�� ���Zt!��]�k�# 愮/�.�v���[e.��{����&�M�c8h�R[�]�Ԉ<#r�{7U����MXlB��Jw?��2�U��@�u�l	��&ψ�&��1/�A�1\'f$3����
�iW4ŪӃ����T�g$�δm��:~��H�) v�4'6���,��R�n�J��2bQ�|'���>0_ހx�si�o��f#�W�N�ـ�A�ѐ
��x��륒��G׮ڎ]lN�/ќ�{i�4�ɚ���Wn��B�I�z���54,B���䧝����d�P�,�8��F*���f�o�c��Ѧ���:&�cy���������<�������6��z"���x'�|E`*����\jSo�gծ���&߯r�vN16S%�6?�P�c�H���Ke���bA���	Bx�~�,��.����6�Fth�~��Z���!���)Y	}cV�L������K��QX�����n��-��R��~���-�XQ��#���9�Ŀ?����hd����^�~�s�M\!�@9����i�q����k���Ï{<����f���4�eUy'������Չ~���_������gP�j��ϯ����k��AWyȬ�t~nǃ�*�8E�����+�Mn�ꉋ�g%H-�]D�gZ��[)�