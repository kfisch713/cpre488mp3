XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����x����Ʋ�"�}OR�CJ�\�}�j*�����i)
�"	E�}��}7�!���c�m4�Z���5���}%��m��6��٣V��x� L;��d�B��*�N\�̔�7��M���H��/V��6���G'������N�QW��).t�[l�
���"�o1�s��@F�489҉�dn�<b�cx�N��o�"l�o2kjDmޞ��	(�XX��C�(FH�M5h��}2�Uf�ιD�e횇��"7�gL��[Ux����>g\j_�5D!�m�ߓ�Z�6�����.?�B�f�|~����K�������J-��l���5O�T�vs��`��3���B<v���(�'�K������1*�O������!a!(���X�*�m��i6��m�D#=$`�H���w�~���RB�3�N!8��,]|4�!lԲ� �<qn&�#x��`�cLA�����=�X��sk��}�L��MO<�������Ix�&H���h�:��Ċr��J�l�ƵΖ
,J��|��2f-L�W����k�5g��;|�/GTm�X�l`��T�w�?��8o�b�b*�#�ޒP9��v�Y�\�����8��6�[MH�rC��̺ꎆ�*6jD��v��}��i$�����XH��T-2�&��4�+�xkY�˸n��n��1PP�գ��<�=��2�bZ
�=�� .�AL�(�:��B]y��.;�I���u|�xXlxVHYEB    1e3a     a20C#�ԐV��P�`��:.g��~���cՎ���J?մ����@S�����
�hΠ�y�E�%���WyՁ���%I|,��`u���yϐ��]K&��>��ޭ�tij��4jS��M���y���3��g��L�4�h��C݅�r�eG�ӿw��j�bn#��"�="ڜ$���b:؂?����@Y��`p����7���\.!8�3�MC��r���6��ո�g�[��M��a�@VQ�ч�$����0H`LK� �忬��z*��Q�N��_I౻���Y@�Kx�^�c�y)������� ��D'k1
�g?(�+ǉ��^�ڃ��R��C3�36BI[�6�c[�)���[�N��(e�D����H2�aX�w����̏�����/�0aP|F=�ب6V��m�m�RI��I��S2�zs;X�*H��XB�i8<�5�p6 81�3-�~�=�+�PR��3YM��(�30�����0�#f5l���sW���OB��1@�O$�Y3���S��ܞ�Ƞ+{��C�_r�Ɛ�'��)��Sxβ���"� �s��b�]�U�36��a��'+�t��w���+�ό��r�C8��.�K�!�;U�{6Q�U�.D��찜�^&)�@_����y�/�휈�n�ޱg��|�]ѣY7se�L�y�MUJ�U����m��hMۛ�"�̕3�����-�,̛,L��fĝ�2�<�9��"��I��G�� 5>5��?Ix�2�8�PecnL�;i�w�a6�V絛}dԆ���,�w+�-^�2��GB>D[�Gj~�ҹ����p�B�;{�ź�!�A(�կ����w�9Bޛ�&�-��bF/!�$ΐ�&�yW?�@��Sz8��/�GoB�8L�RWvF��qRP���BN���V��W}�3��ޤ�/�.�/�_(z ��Pcn�q����+�`ک�2�VI����$��9��&��$�3�S)7�^pmU�D�S?Ym����f�������R���4�s��|���\>�I�m���t�82�,U����[8�!jG����YI�-(F��da�%����i%��r뷂t/.%�0!�ɴ�Y�r�zh�"4E4�Y��Xk&R(���؀�⏉����/�b�x�]#�)#���U� e�U&�ۄ-��SBmW	�Y�� +�BKd�A�����w<ػV��L|kC���W���/Ԯ���b��ro �{ٞ�q�|)H'���<��e��)�*S�ff�-f@에��4�V�b%�$"~��&7������P�t?�!9�	�q�& �8�+�[��xH&-��Ѥ�٤Vaۺ_�>�ʙ�ދlGGV���66A#��{8T��2�%M�xq���4�u%6OP.lx2� RU�³�3�Q����)�Z5O���̠p�
�f�
�	Ot>��6?��x�&�0��)~�=��{c��R����U.��E��[&qu��2���$&H޺���o��%_���?w�'|k�%g6Q��!�HL�T�$�ӏ��\GSGx�_'p���`+^o;Yf�~
�!)O���Potȋf̸���+N�u�0�+�j�/g�7�vn/�ߎ���gN��t�`���&RF�l(P��f2�{����5���Z��rTxI1��N���Kf�A��,���l� �1WL-���aRH�U�S�[�=�Ϝ﹧In:�I0s�F�:MBh�WjV���֨i:h�؃� dE���*�\��)"L3Q��PyP��qe�nush�5�3���s��^�؃�7�+���<'�9.F��`&-�C]S����:���5$��;HG�ґ?�v���{� �E����1��!},h|�{޿R0,�Qӹlt�[���ڱZ��{*��A{�b��R��lR.m�"ԣƠ=��O���2��<`t����繭�|�=�J�B�n
�*[��.d[e�������8��X��WpSO(ŘU�����}�EL�������<�^ �����ug�b��]�W�� ��-İY� 	��4��8`?��5p�B����'¡�C�2E>~@�hL�3b�4'ۮ���ʁ��!���J�5����B׸T��쯏j�1ӧ}Ou����7����G
�e�]�Wڻ��B��;j`7���h��N���� �m��o��1l�b��[�l���!������	
 ��E����q3�`���WYlґ"�Rv���>��D����S�R�M{BN� �"?���6��3��<�fV�!0�1�4��o0��D���M�p�־�g�to=խf��B��b�#�v��9�rb�J�	�����u�[�E�X��`tw����x�@RZä��m�5z\ꋱ��y%{��=_	*(���p�Em�ž��;	⤾��מA8$ͼNR(X	��q��S$��3r���ݢ%Oc̑O��wu��?��B��j�*He�Qxb`Ӝ���9�ʘ�t-oҝ�?���Re�CL6�٥C��� ���&���	"�4�
�0�{�5�7?pX�-��a��<wh��>��-9H�k�Ʉzch��E