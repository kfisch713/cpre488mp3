XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��/+����CǮG U�~��5R��ߔ�i!S�q�={A'L�F���N�Q`����v�T�j��2=�u��Y�Ϋ���/�	��n���!)W��eUL����뇃(�Wr��.A�iF�a����h��G�2 ��i6�2���R���Z~�]\�j�D��%%|��l�����m�8���ߚ�TK�������B���
9��H����������ݮM�4~Gt���U%�6��Q}^^k��Q��c��TKFC�Q��i��TA�K82��5�L��yoN��Q�R��Ԭ�xM7p�'\J��f�!��y=�2bTe�, [q��X���X��/�dr��?Lr�l}ȴ�ҿ���4��е� ���JB�ׁ�-7� �������p��� d�G,����4n.�?u���7B��S���l�TÛ�Ǭ""u�e�!$��t��(K��¬�!C�1EO=p�0�e������bY��ކ"����-#�
��;�cD$�3��˞f��9R��{��FR.0���`h���=��
�}aW��]�aV�C�X^on���ƙX(�����k�&m���So������Y5�]0:�*U�kݟ��d+�m��`��}���a��][�%df����]����@�-RW���Ip
p�ıѳtp��Kp�X?���h�	B��4�C�ɛ:Ʋ9|�K�:����v���pnL���{�Ȩ�Z)�&�'� �|_�P�z�b�zXlxVHYEB    1847     900�t�.>�V�`�V�w�B�c�H�܀�l�����d3��m���?L��ʜ�Zg��7�_��/̙���+�tfz����O��(kI�,򦜙�$`�E�f�x?�����QS�N�f�c��P�0׶�Vϧ��Q������᯼	���N�+��V'Yk�E1���آ41�B���>��x��:Y{t�1Fm��e�-���8��unO�<6����K��	��-<7�)�x� �a��h��^T��č���C�'.�rN�k6}1�:N�F$DQ_�i��Ԫ�4.A2Sl~���\N<����,(��Y�@��
�f�In5s���T�E���>���y����wZ |�F�8J�p|czҕm�3=w4�`G5��1��tف&]� �w\S�e��,�F0���]C�A����7j�q' �P�0�`�,����]%j[>no�=��'z��I���$!�.��zF��,S����~��d���*���*cT�H��(������-�lA�2o���V��+5��Q�O�E kD�2��r���D�n$$i,����$T<�s��#޺Z��-���� �a�P=��p�k�� ��5S�>ɍ��a^�F?��ߘ{?D�~U^�R3��Ȋ0	>TK�����G�qJ-o�m8)~��g'�-kSK�"!�:�MV=������m��!�]�/j��K�B�lI��0�q��%�a�$;���5�')��V�[ &��!><�&^��\���U����I�B�o���5�=G�a5�(�����b*�UH���(ڭwme��)�21t��bT�?E�/�ʍ^�SsnN-�z�)O��a���%�3%M�c����Tς|��c��E�"�zf�*q�<O��Rx������іVd$������F�JB���e�B�������r���؁cBۢď�����[Br�i���^,W��ư�f�ڜ�
P4�����%�=Q��6S��*?{[m��X�w�z���2Z���ں�t�b�3Mu� o�CЃ�`�:{�)�m��4w�Pͭc G��gL�_�G`�*Aiŭ�������y����Ů�Φ���"�����ӆ:��G㉌x5��-�SX#�DOx�=Jr>�Q�,�������S�)���Q+���R00m�5����\�H��y/��#���+@0�R�wu#���X쌻,f�n���V���f�����p�3}rC��=#���;�I��\���`�K!���򦣇�����q�sCS�A��� �""�?sϴq�>�)�d��ß��7x�&~OY����x)!14xE%���E~�P��+�X9'#��Gf{q��A2����Y��l�����`v��Z	M1��Ѱ���"��1& о�B�)Ԭ���k��磤=s���t_5���ED��`�	��'�hW��>O���%����s���S�H��V>���{��.R�":��R��9����GX�O*|�Tq��� �Q�p�ʭ�;�X`�_#�������활d|�v
�#��f6i�*�}o1�|+%���<�QT�K9EQ���?D��ID]�.�:ׇbT?:�#�!��Н7��,�DB8yĤ�M5?�
��~�m���X��\�ڦ�h������>c{�3�%�d��98j�*=^,�|�|�f#�Y\��ȷ���6T�Zq�8�֌���H�.�plfya�L�p�B���$P��'��}Q���34�l��E�w��D�i�3��`o�)����>;����k�&�*�~ȡp�����3��yv����H�.a�6>*<8���	<(s�â�Y��5(�">`dv���b�v;����$��+��{Q䲢ɑݹp�� ^K�7%A\߆#Uj��q���Z@K������"��b���R�D�PJ0���~����fZ�l�x��K����ν��i����E���<X&YV3������-~�0c�{:P�B���_tF������L��%�3kTz��''�F���j6}he`����j;ժe�3{q�İ�m$H��Fa&6�@�:tR�����~�.6���o3�����+S�3H�]�&Ov�ꁊ5�h��/7��F��'��iG��R�*IN�
"1z 4U$�X�[ ��<>zK���ئ�aZA���l;�f`r���I�K�����s�`N�Ikr�
?p� ц# j���%#*v��H���1�8s�L��Ow5R'�f���yw��G{%�D7�>��<�V��6�U��:�[�2K�,�H\��