XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd������CЍ3�QA�=\����I�A!0�:�C���g�3K��-���:�cT ��^D���;g���	�����G�[_���{�[����i[�	�pm-:�~ת�����G y򔅒����jc��������z�ɿj��h7ߢ�:6���I@����R��������ƿmό���!W[�)~�"�9Y���@6Qq>ǡmI�$<��>#���s�^4F1�X�iZ�?���x�<�K��?$�`������Ғ�Hg�������Ȉ��+ H�g6�x��T*D�Sa���G����pc�y�d9�G��_`��y;=$��c
䠵����Dw߆,,�SL��m܅p�4oy2��1}��_Aڋ`�b�_RT\ �:��x�b�!��KG~й�5��7=mGHG����X��#��((ǡ��xʌ� ` ��P��ė2�
H��kG��A�u5�؄���	�C�d\Vľ�/���$P�u�tY9]�~��:ϲZK�����ْ�[0#�ٯ,<�SE�����.� �]wѬA=㾞:�/%��ktN��4H^}.���Cjb_�ǆC�j�n�m�`x�[�.������^#��%�12���@�P���͓ţ�_�%0��(]��(�B�G�D@�HM�F��uo!Uk��r�"iy=|���� m�ȸ����c/J!-(��0�&i+��HÁ[ �L��l�"��UET'���+���a$�Ɵ���~�-�M>�Lb��Z+�J$P���C$}~��$�k���ZXXlxVHYEB    da59    2e30U�~��j25����w���]\��.a�h����C?���^��^�@$h�1��.�����j��<@1|��`qN�!H߹>�k%Ȑ�k���/}T�>�Q�&���ҽ��w܇Ά�\��J{ق��;�h��(�2W��?{�n��Wr1'��1�KO�8{�/o�\pZ*�<�ѥT�����|c1��:��FM
N��Y�h�IPų���7�\��Mn��z�l��,݌�@%c�uw��� ���a�=�-�P��0��f��+B%�?�Ň�Q�ր뎷����]����ܤ(E��R��Ku���ƈ�F�˻���s*�H hTS�����b�b������:�5�┓�w3� |�5�����'��C!��h�A��(�b@B�GR�����zY%���]��W8jm^V��<��6�ƶ��I�K-,�7yei�����8�ܠ{�A����=��i�-��ڞ9SY���>�ઃ���Zq�⊻Lc�R�H��E�����|x{����d��F��7<�O��r/"zFQ*��O����݄2sw�v֓ۨ�B���n�����j
w���ҲC��4��R���د\M�kKK�os�y`�ÿǀ��n)�F�R�A�0�I�2�8ېcq��������kwW8������� ZGſؔ��̉Yw������	Q
�(��O-��$!�x��(6!�cب␐�I΀Z��{Am��+`1�9�����m�@��%S92�}�|�bı>��U{�͗�3P��=��$%`"��ͼ�pv�	�J%N���0�J���
����������LWLT�|�>n?gQ(V2Ԏ�r8�<D��V@�x���8��4[��O��?C(rL��!���;":�����?t �|W3P��UR�L��~�V��z�h]���@C_�ʟ-���ԆxQ�����t\l�M��|4* ���0N������r��XN��@a��������6��-�΂T�&Ae`��Ւ�M򜩔7��RF��_����Py�}��k,x=wQ'�n�uY v�,Q:C�rp�����K���P�9s�ER��
!�<��B��4ب�A�<I��4��j�;��R4���J��{NgA�UͫQU�/v+ ��HFcc	ֿ�9�1�ت=1��FV�&]���E	gٍU�Kᷖ��qp���)��(u�]�z�٢�/��(y/��7Z�>����֧0@��S+���F=�e=Bx�{�(H�;3���asw~
��z�"l"#��1�Ɩ}�n;�;Ҟ
ND���Rv�s~�cB�%@��RZ���w�^�����	yx��)�d�a�dF�l:�i|�Jp��.k邘l]� b�`�G�R{=�Й�Ei�C@t ��l`��W����5l��yO�*����X4Tr �K\=��OzT'��%-+W�b̏5��P�1�:�x�����<�����=�¢��He �:��2���F*�K�� ��a~հ߾^�S�Juܮ�?g�Ά�2N�H6�n�M��5���ނ��/��+��ҕ��&?�;��s*�M[�P2�,���������=C�쟇T��2�	2���7�2�2kG�F�}:�x_!��u���)7�I�k�x^�/��{{��wV�C=mx'���|?�}�3#�_�@}�섧#�'�5�k��+���O����{ ��X��!��-C���#��i"�J;���F4,�m��Z�vF����^㌭vqy�1����؉�GKCl�3���r1��4�w��Iei:����ey�d��uT
���xt\��wDD�$�C"���=Ovi��vKY����l�s��D����C�ذF�[7�5�˂�����/;�<�� &ʹ���&�F�DUu|�4�p�������w��o����w����b���g��y�L����C�ﺪ�p
�Y>�ec�*���V�7��p�P�h �؁ǀ�������*h4��/�=X���BIgkj�l���a�f��S����CͰ/p|^�#���^��TCx���ye>*����2���΋���C����kgch�)�6�A��&���!�1^��|�0�ٻ2{�H���Zy����~�#��O�@P�����ԎtK�-7��OKEoz3�lG9�Iz�!0��Y���b*��܁*�/{���/�S6)��[���x�lf�xp������dض��Ae��b���d!�j�*��4-5��v�_Cz��ʌ��y�6]v�V���o�`~J�@�4���m�DƊg���.��,<:"@)��إ���s&  |z5:�q�zT������u����8�I�d jnh�;m��9r�c���9@O�|�۝|��o�A�Z[�d��3����+�7�7I�TE�kX{z3}01�Ӡ�9��r�!\�G�ɕ��A�k۽e��w`9�yAqu�P�B�	.k����щ�X*w#ɒ���Ƨ�q3��uot}��,d�������1ʭ[,����M�v�r���]��	*�����&1#���S���6���r�Ui�,ԭXx:�!f2ö���Mf'�0z�#��|{I�M��W��5K/W�T%�%ȕ��Ԛb�)�5͑K���±�#����Ľ~�r��Dj�uj���(~t/��}�/�E�(9��;���ҭ�}W`��I��D��cZH�����(d��K��
:�Ӱl�f�FB��nI�*��)7�'{�/wɻGf�*�Ǫ�-T��r �``o_�틭�or�VE��P��ϛ�=i���V��FB�l)�h���y?e�)!�O�f����U�9����nʀ\����ӫ�V���z��� X�F�Kk��z�n����Z�ka7@�m3�� �%I����9��aI�)ur=5~Eg�Cθ :�!k� ��Ð��p��Ӎl�I9)A�؎����Hh�2�� �/#�`��1�mq.��q��E L�J��T���N@p�@��}%�S4�ҙ�gװ橈&��B<vSV}�[F����u��`�31�ܠ�#DB�Ѽ��S�9pO��8��z#E'��g��?�n���g�XqBO�]�1��.��!��[��kZR�5��?I�B!:-��Ǹx��%��AF2��Y<^NIP�i��C�W
�U�����ŉⷨ���N�jf�(~wOb�+����e���(��������?���yl�F,��������P���}��L�!�3�̫ZS+�c�������\�>G���K�Q&It �`CF9��X�s�]�����|~����P`(��BB�v�t�oHCWD��D B�G��c�!�{����Węsp�7Ȃ��7�$_�5�`-�'�N�s@j98� +B#mL��E�>)�9%S-��� ͂���T��̃�+��V���&�Z��P��~t?9L#���D;%�W��x̔V.;�=�����-��Y��·|�3wk�rI�|	��2�5o�$�8sX�{ُ���؞|�� ���h�GN�:)#�����nl����5��Q�<��g�+����1a��	n�Œ��Ov�>b-���z�����B���XU���VAx��(�����8�m�nq��6e�7�u�r:v���O��s�Aګ�t�\p?t���uE���WA����X��8�1�F7l<7-j�Yw���g�%����Ov7�9�z�L��-�c��O��z�X�Hn(�4Y�:���' ����4(3s�Y/�x����:"����V�W�3�K�ҧ�y��Ƙȥ��k!^�5�8�x�"��C�c�MkĊ�;5�5e���>^4O�U?��3������,KR�4�5:
�1"5c��9��Ў�|`�do�Q��r�l�c@��0jɤE��)���4���?q�0��IN`1T�.g�O�o!,�?N���xҨܜ۽�=�[��0���=��d
�x��Y�nhZ�"�nzu��q>�C�NY�>�【>���G��g6yJmi��n=1�9���!iy���ñj�̚��6��n�f�hRj�"�R�m��f���h�X.d�N��Z3�Y~��J��P�	ou�RB��W��;ŕ`�P����O���f�b�z���\��+s���+��Ա�=���n���׻�R�+^��csOS���k4�kv�c ��˼;\e�dU��_5b?J|A�~���j�!�����Yԇ���C'�⮉��K�ͫw\@�	�ƨ���Oie����e��~���P��X�a����k�E��@�=;
6�ߍek %;��v��wm'�C�*)؏(�d]��f���\YƖA��l���Ytg�n:+���W0�m�y�f�>0k-HP �x1�t�)'i�TP�-����~S??�H�����/��B�==����&
~����ëݔE�<Ms�ss��$/���Rc\�'��Hw�0K�u=c���J�IU����/�Tc�R�hv:��&��|y�jM�9��ʪ���cx'���ӳ{�bW	��hQ3���%{|-2�C�R�(�Ĳ�@@iW����F9M�o��'4֕�%�u��C4yΐ�?��ޖ�;!���=f�쒲�=��}V�p����B�h�1$�U�U"`N�5��(�H�r�q)��w�M.�@d��A^ydɛZ�l<a+�@4�x�nM�X�ˎ�2΁�c�B���ܧkk�j.��m�VD��_����[�D��EN4�p�R�I������9�%���1Hb�l�.��,��}G6Ԏ|ҝ����U�偩?��ݐ%�C�<8e@j��.��&7{�5����(j �߼�����9��Qz~t#�ćdM��r^%�I3O�%�:]o��W�<N-n���U va�|^�H|pi�����<��&�G6���}i��\��e�=Ѷ𯅵��;�EΥq��	�h�ҧ�^;c�ګ����ϱ>�P2#2�j�c��
����b7���� ��+�QD���
A��D΋�[�,YG�����A~>^�� ��*�-�7���
���u�Z}ݾ�v=W]�$k,�GH�,u��0��	QZ\�*:��T�=T�Y��?+�b�<a^��F��oMWqBqM�GO�%�1�c�u���pv&đ	�Y�(&W^�R�u��S�4�o��~/ �3�M������l���.�(�e�kV<�a��eN�]R���S������~���I^Z���Tx"�/���̬m^�?���o����W���@Y��s["#�B.�|]��|�����B>� ;jqo h�8��S2@�WC3E��$o`����׶E��0(�^cNH���2w��ɟ�n�?��\�מ��y�]����H���O���e��Qa�+�#/�E�rc}���B7/��X�����G��zi@�9sY�P˻�jC��o;|'�y���T�og�F�z��� 0<�4��\�L�o B��N��'U����*uU�@u<��=B?Ӫ�f��[��Ȇ��xȞ%��Sb����"��A�q���M3v"4�u��O$��N��ܨ���,/�B�4����a$NU���x����6_Z4�2FJn���$�"s3ӗ��u?U\�~�c��m��`�軆!fb��ր��#��ŗ��%RHZ���x���G��"�P��nYsWaI0�r�r��"`�� y�ޢব���_4�z�B�����:'=H�*������4����m��������Ǎf�r�y�)ߓ��dd'˘�L�w�|Y��V�����s�V��%9�5WŋA!�k��oHo�-��Mq=a/�k�B�6✴6�a\��ĵG׎
��%����җ0��f?}j��~��4��S"[�C=P]���6��G�O/]��Ic̚��`�	�a��!Ѩӊ�}�\�Hk�h\JփUM��QJ������>�����*�3���G� �7'��-O�Y� OL� @�!� A~�2�9�H]����:��̿j:jBY#�&�3$���,�P�&��7��&�5��* �P؞���Rʘ#?(_/F ���� ��_\y��~�t	� F,��hzSȥ��Y�O�Ż,j	1D:z�ԲW���#o���V���0��|n���U�m@<G�0�֥8�'4W�@�M#�z������Ta��'k�y⾣�͙�.rĻHZP��]
��LH:�a"�5��y2K�V�F}�����;޸�>Û�Z�^Ө��+�q��І['ҋrI�l�9�;FH�%�� �)�X� XuPx�ua�J��Z�ʖ��p��e�p�_���$�[=jeM꯽��J�����߷.$�i<���@G�~Z�$��&ö�J�����*85��X�� Ps+�Q�w {sn����X
%�C�*�`�F�����4�P��k�
��6dc*�	�=ܼj%����P���4G��z2	@ڔ'�J��؏�>��)���x���n�*�p_G~��U{h	�`I����Yk�,3�퍥��e.�׋��z��[G�!��	�f�o,Y�w�<�s�QQ�^�)�+��uU�:���x�@Ą�^{yB)s��='�η�,��V8�J�����	�)X��#��S~�DlF����x�Ӛ`׿�	�>
�3"=�/e�.K�d�E���M����Ȟ�k�i<瞴��|4��#x�HK�4-7����b��y�/�ŭ΀�nY���;g.'I���O[�W6��ûx,[-&D�BjW8�o�6}j����z&X���E��ȈJ#b'>ʨv�i�9�?��&U�ke� ��$�|�ڑ���X�9���88�B� w��`~�['m�_,�����d��J�� �@�8�v���lY�����y��El�jL��i)@n�G�S��A '[�-����^�ܑ)���\�3�~3��l��iK�%	U�vDȿ��Z�|���nHå��%����z���y=G�`zs���/�P�� �&�A��&Gyc��W�nӵ���^z
�	!�km�[|y�a��&�n�p<Y��˨m'�C�qG���Aw���qX
Lt�6�a޻���]�C���;a��$H��G!�݁��s9{Q~66���z0i���'3��;ǳ�u ���l�m��vw�2��a0Ql8<¬#L�:�Kw�ͻ1כ</=�TX��8���.��H�WAQJpp���!:�O�Qƒ�G�����������S�ț���|�z��	q�Y=5�������T_���`;6 �)
o�̩Ŭ�ڌ��Ƭ�r�v�l�a���+��RmN3$���F�+��g���:������E�nX;�Yq`и�$O��zQ�����F0�(�Q�˳��Gp�0&L�P���ƛŊ�	�8�������Ak�p�۪Ct6A�_H���q��+������)������q&W�.)�4��0q�v��c�񟮤�����?ւI����vl5nM�-�zk��v��;���{�H�Xi����f�[����4���{n҆�d��Z!>��E �VQ."U՛P�CI;��WKX��pLy��l�� WMʓ\��Zz�:�*�V%k�e*@G|K��ܿi��J��O�Q��XB�����H*M�ZsX#޿�n�0>��J^�g��p�r��>��)d��A�y��d�冱�MnX�Ds�����_�0�<4.�I�㺭��3ʺrԈ|�C�@@Y�«7Ύ�?��!J9Y��!���Zv&��c�Wt=�5,wϘo��F!��#��|�����~������hP��s�m�R	:���)�� ����e�XN�JȄ�W)�ۜJ�Y���:Ĝ��a���Gܗ啞���ȿ^�pÏ��T��W2Jrr��9�~��4�5ԅ�,>R�J�"@VMwW[#�U�O��??�Ҏ��þ��
����K�T5y����?.p�C麲*p�P�z����ys�_-#�_O�Mqz}��?�9�,�D��_��W��\��<�a1�4%��j�'�I��W�SS�sG�3#YP'��9��P���b�V������I`�y~���QW۟������y�v���!'�e�����s}�!A���7�۸k0Zl����qʸ�.�<��/�ț���T��Ä�5�I�w��N@F3 >4J���`���A��Ω�0�Аzʲ^Zq-����-������Ő��+�9�����C_�P� �
�����an��["k�")
�D��=Z�O!g�HM�o'𗿕�BO�1R�ZE���8��D�t5uFA�����pEC�O�Y^��m���@�0���?���,��S^�b�ܒaQ��_��6���F��LI�:�!��z�:�ڦ���c����ȧ�����f�S�<�Y۟2�B��͋Sd-X�hۏ	��ސ��f�W�C�x��J�8�[A��V�]齊�)��]P?i�r��U�Ы�$�� �p��׼��"ՂW����۬������X��۳�'���-��_�����]�B��c=0�4�YH�b�Mi��^#�)��c'���}GvK��Ț������'$d�UA�=�$��_�p��Y'K�c�A��HN�=���(}����R�:B� A���%��'���È������Kb"�jv騖�mr?�;�7JW��Q5f�B�����+�^����|�4.�6!��>(��W8�����P'xB�8����'�?��g�$�� ��eO����s��|���C�2drn���7�����%2Ev��Bw@Q�#�Ę�QC�YD$�aT����ǹraT:���#:��dqh�@3���B�B�>Oއ��Kc��DA�]E)#�Ҋ�Z�ǟen�F7��P�[Ѱ`��q[7kܹ��U✱T�����|�'�	��J���>Y=V�C���P��A�Q$��hh��=f�d�v{A�`9�L��#�k���� �Ţ$��1d�v�8�. �
c%��g�*wf������߽�&��H��#���̖s�j!�#��(�A$�X.�O�\�A�HkG��)�'�S����͞�Hb�{��M3�s��\�{$�Y�̝���p�Z����,?����
��a�W3�Y�\32��jn%?��y�^��1�(a$(ai�E#Ak�8,f!:�T�	�v⩿��M��S�æA>O9�^{�_f�}�� ��e55]a?69�1i��Y;T+�6�+�^�UHf�E-)5��0��i6�x$��i�Hą>�w�f,;c�����~f(�(�b�a/zEl���X<�����v��@�.gE�lo���-{���uВ���Yf6Sfǀ�Ka��T�=-�P��~j�����PzS�|�}���e�ʱi��eA��I� �<�p5�:��fR 8>x��;Ä�
��S�S�;ami2�@�ʍr1Q���0�E�ۃ�y���Ӻ��nº�&�4_�c�|RL��	6dp�L?��l�@x�.��V��j����#�u�"���@��u�����@�n�:�Ѥ�!�W�<��������>+��k�6�m�k�]��=!�[���3��	#Ҧ]աupBX���'�>�(��t��R��/�0=ʗ�#���̐����;:ӝ6,��t�1��>v%�24�$C���:�x�k���@�v�*��{ob΋}'1��U_� �[�~J�l��z;FCHǳ>.��"���ء�}���{'k����El���G�CZ��G��_�Y!��Xd�=V�����5��h�hsS�F3�g#��|ֶ��c[�f�>r�Jlڌ�4����8�|�.���r�uac�XhD�� O��LP�n@��������O���=�z,C:O\\�m1��)�<��[O܆��S�<G���'X��W0��l|hș�HM�qc��j�-1Q�Ai�`,t��⚭2�Gc �B��ׇB�v���Y[��pD���UN���rI��T;�<�[!&��Fuz�]��}��1����)a���G��p<�g��K�v��4��רGmB%��\�b�n��ž.�_�<����.�I�7�hf9�<�������g�Bl.�#�$�L�,*��</J���>�#�H�o ���� ���9A	���Վ�tIܪ8E9���Yi�;3k6�s\�w�ljUY��r�dѫ���y�|���+Jm=�������X4\m�ʈ��W9�x����9�����]M��<y��MF=���",]gڦ�>��h�� �"s���	x�)�VT��T��4����J�	1�I�woޠ�ӏNA�l�eCzVzJ�Pl�]}a-�����'��\$˷�f����}���G��Wimʖ��A�oW-҃Ѭ���;B��)���{d�|:=%Ep
4�k}�px��Ne����楲%d�Bp�NJB5�|ن���@v,�Em��P2�&f�^�Rz�D��V�]?�t���2���9��z��7���M��l�)u�5�:�(���~�i�$VmXi��:�7r]���&����eN�r$ΊE��ɬ։��@EN1�~jT�Ћb`WT�y�DG?���v!�@��0�(	��D�шh1pK�qn�o�<su�|��+_�q����>-����� D)O�[����B`j��dd�j��_��@���Y�閛rG9�9�wF�jZDU���uMoi�BY{c}���W��z������� ��$����Q����b�I	�
~��p���
}�w�s�qu�>]xn����g.��gx��t��zI�sާ~F<W ���ae�lF�Ra� ��zЈ��I�-�6�_�=ۋ�Fb�6%�♣���@�l��͐����q��:g��)\�U6;�<�5s��&f=��ji<�+��(�
�_WAzA�T���K�Ρ�^zp����	5�a}�s�[�/��o�/��T>W�u;Ņ�v����b�S���ܹ-�d�a�uB�x�tI�7e��N�M ��.�Ĉ�AK�CZ�J�Ջ�F
Z<�dTE�?��K@�كv��`F��hj���=�v+�O�ئ�:���}��G尽l�:_%e��y�6V���w��?���4-�Bf�i�P�Xٙ�%($�z����3󶄆��������F3�{���7��:���~�)���&^F��`�`(�L��*6(���"l]�̌���ͽ�*�Ý��ڞ�&?��-f�³�.F��ۦ�NRi\t�!.�H�ua��g�����o)u�C�e>�|�oX��p�R�����.��$&�^7�|N8�w�����b�Db���ڱ����n��-�-��]�XuL�5]�V5v�����4@]�	�Q �u��D��Z�`7��O��j_ԏ���l���|TK@��L���-��R�~���0`�vG��o)���-al�����E6�v�Dj��p�����Ȭ��z쥕���|6�Q٢��>���b�p�~J��?�����_[̈�h��ydI�
eӡ�ё\*� n�#i��Xo�4^�+J!����X��&JX:�$�?��݄�3�,'�$�mē�S3�j�v�{���9H��"$��&����I��g�.�q�.G����5]�����8B"�>��hF ��L��Ir�x��.Qiʇ*=W������{	� tz���A$]Zv�z��Ų�o���=���Nد�kU���i�E���б�F�}����=��臎�BYǃ-�#�'V�^���O������8iKujg��H����{,����(.
�-ѱL�O!�C9���4KJ?C*.��-�k���R�P�س?