XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��k�.��l��%�zY�PR�V�\+ݿ����
S�Ǡ�S}�֧rs�n�\��Ƅ:		���//tTI��������?������Rt�{�N	M�'�b��{d�KU9|,��a��	�W�:�2�l�t���]r�~d�9�쿓݆ r�ӦW�,�������z��כhT����_���혜�`i&G�oF�T�ų�(�<�l}w�-w��i�$�����s����o��u��fGH��?ϊ�=ޛ�7&?A�Tr�q��))Ę��Qi���u��5�E�OR]�$p��A�������gUfT�Ϧ�Z�8ӽHz�4��r��;�<�j�a�%U#�C���Ō�c{�bv�+�&�زE�}&a������R��M�π>�ۈ�|�[;�\�^84��eU���4�x�F�/t����"��S���I"�h��9�ju�A�؉�����F���m���S.��x�h�i���?� g�\"�VE����_\��)�z�B-�C��w.�U���)��B��#����n额���ؖ�:{�,B�&�uUڌIh����(�~H#����[B&6�)5��L 5�˿-�"��wÞs�[Q����H�q�F���ifAx�Cƾ�=/|�^[�FӺ�J�D-���X��J�txqM@FV��q.��p5�]U�����As����b��S����\=�%qP ���K�����,K>$�L�q�G���<~�����9#g��V�
��-XlxVHYEB    3b09     f80�0S賧�1}�d�VР��5o3Mߧw��#f"�O�tf&]Cq�*L$#����{�	v�LγAL�mf{��9k�B��e�Bqw��7�6�Fh��#[/�ՀНFmH��0�P�g�u���O�]i�D#:��g�1A��
<�Dzf"��Z�������ç��N �L�"��+���vy4��(�[ᔋ����_���T��V�.Ż~�k���}5���!��sw=Βʸ��FA���S���GvA�9��.�f�<א�|TKV�`I�4�:��<50e[ȭ�h�V00�
N7�$�:�2Є0q�F�\\v�@Qn�٫����>�26��n�o.���:^�����ޝ<KOpi�O���W��p��.�� ����k�XdwG��R1Z3E_���:�nq�mIL�D\���C̬�>`H[�_;���QA�/RV�FQ*�Hq�H�mY���FS�����3Ht�Q��\m�Đ�j�:�'�
��Ƚ�"H��ג������@�?3��&�\W�!]s��s|�͡�E���gwdb<Q3�RV��_H���3"5&����H]��8�T���^�q����*G���PAű%.u�1q��-�p��oWGiq��>6��pp��^���������qL��q�nŘζ:l�hے `x��(�z@\,�|��ډl�������R��ٽ�v�`h�u���@�pݦ&F�����-s�I`��"�<���x��%����غ�P�;z���Yյ|�SU�Qf]3�gs�>aS�>���Q����-9��?���3u:וؖ�0xR�n2�
�� ������1l[�)�Ο�rC}� 
7�d�p�zW�(h����)-��٠FF�_HU����%K��X�㾅}w({��Π���P�9[�����jG�q��HZ:P(�������V������a��N��p�t�_��~h��t��J�M4�~]`�hи��ף�lŋw*gCCvY�RL �������gإbvrX�H�U6�bב
(�Uy������򉑔Y��Z�3�	�P'DT��̏�I]����� NzpZ��L04aHC�,pW&R�T[�:?��v�^0m鈨�����fگj|K˼9��:hSv�ib��֞��fK�	��Ff�������w���Ge�P��Ԓg`; ��$
d꿋�&~u��ks{������ux^$e�e��AsqI�X����+׬"�[m�>�6W�;��UR�ƃ:�U�@�fa��=��zYCR�^�w%:�DxG�}[�>®I�x���T��j`���un����>(�I}x|�x��q#x��_��9~���B���}�EY��;���_��Vu�|�ؔ�0d��w�r#ɗ������@Fx
��W	�k�Ɨb��=R��̃�s�:��G4�A	�Ox�:7E�Z�v�:͸G��CI���R�c8߀�eB3P�[{�䄀�0w#��TAxM)s��P�ՊJt���"��?s�sm�2��� �K;���nq��T�$}�7v�EG�w-��8c�u���n��.i����Vz\��LR [&�D���ѯ{�o�`��gzj4�3���n=9����ip��ծ,��t�S�&(�5H�_�7IUe��%�¦L�PH#�].��b�-J������i��:��qQ��W��}F�Բ���.�{V*]23(�uF��O�XqL���^@�s��Z *x��ڒS"��̬�$��A���\��o"V� %Q�;=D��	Տ��8�N�@`&5�r��&C��� �B6s5HN.��������	\�+8֙�IEa���S�!���-��L��=��Ŋ�4�	6�SӍ�;������+NHA���S�i=�ͱ_}{B���f@;}�D��3Tg��w
��KD��[�����x���`��D�L�/d��Ϙ^u�pJك8F�HP�FY�"�Ѹ�JE������]t���{F#�1�sQ��W��7:I#�q����3s�c�Mh�gMtN���?#���d>��t�T5a�	�S6j,�UƄ�DP9O�f���>,���w-kg�H����ٔ~y�u��"T�A�&�$�n��w����&&�v��h(��6�R�c21h�ZI��ӢU���h�;V@�E7Q6�+�*�`M�Ö6=�x�-��1�8N�H�x!���fH�ͳ��s�l)�ޣ�����H,JZ!uؓ);OZ���@��P4��QJ��Á��؏���H�v�.��!眈����nk�aKT���䓓8�A~mb��Z*{�q�I�җ��p���Z��qDEgP�B��У��>��7;�rt.TPi�E��,�
q ��)���/���Mdct;e�}zrJp���me��lAMj�:��6���>�V�Zq>ь�P�_��:���`�%ߦ&��˩�:�~4y���(�Y��K�d[��峻mB�<�k������i���3�z����ؔmĸ���*�:`�D(�ܕ�הx���	��)�Vr&��Y᧙g>���q/}��g���8X���6�z)MT��U�J�P��A�"�^�:��m澳��q�+�	�P�u���4��=A���m� �ϩ(��E�wu]MĢ#�켙O%�MDw
$�S6�J�5�$������6�&|u�x�<Ho�4A�Q�g��m��[v}
�	L6ŋk�Ϳb�k6�:��bL��5��۰�6���~�D��6����	)F��6R�����u%�f�]��*�BkYj����p�IE%�$1��ۼ6���O�j
�(i��U�q�e?t��D߯�̑�s���oӀ߄gމ�16��*�S+�Q�'�R���y�Ȍ�����	V��
�V��ul'ا�f��+�/��a@]%�;��4J!��.�.���M�}�rގ�-g�l���?c��G�d����(w�ѯ��v��!�r���l�~������T���糺3>�H������U��Q��?��A��qt�-/�b��k9Y<~2}��֤%󐜇�Ƿ�i��Ny��BB�=>��9����:�쾵J����o	�>�ǿ���������gO������_A�)��s���.�.y}C���6���r<�/��p����B��Ԕz��gG��?j�^!�<I]�ȋ����!=T6�U_����#?s���u/%KbfB���_9���%F?�<�A%6ձ�cj�=�mv����gehMM��ҿ1��]k���\23<��|��]����D�Aԝ�H�ć!�ڼ#isrƝM��ف�	:2cX o�?�W��t��_�����d+}��_�M�v�@�
7�fj ��噫�42�m��|U�u�œ���'K�G��ݛJ��,�S\Ks�)L��Pq�ƥ �=��-�2)(�o,����� �ۊzqkY'�"�_�P;�YJ��\�,�VW��4~T98�ȣJ ʠ�}��1\��� �K����������'� ����_#a@��~��Y,�݈�B�x�6Nd�:�w=�y�s
�����;�L��(TE����E0<Qg�aW���u
k�l�w�4�_c��в�l_�v�3'/�.���+;�wŠ-#=C'@i���y�	�fl��ކ����|�jeL�P��u�~�7"�?|
Y!~r �[~��4,X��"��+i���q�s/��ؼ(#Vf��L졔t�x:�I�m�%7߆��sCʍ�=�*��hUE�U>�ԣ �H��7Z�G^�;8G�}���&>��B;��}� ɑ*v/�02;(5�{S ����LY�0$ޙʪ����F�nYj���%�_8���y�B*���%��Q1�61��3��1��MG׾{��׀ЈHpx#)��A��lQ}�H���~���o���]��n@��㏠v��29��M�i�o ��]�`�WɕԨ���4����l~���E����!�.�Uq�+"����c