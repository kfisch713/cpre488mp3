XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��0QQR�l��l�°Ā�۠�cD�*�M�.��&�J�&�$"���/㚀K��������������X��Xs(<����!��h�&n��	��VO_uL�n��(�L�8F�.�[�-ڌ���h�X�R�R7�����:��*���z��7ޡۘ�Cq�IͰќ�+1[�P<��bHr�h���+X�!-�r>�&q^,J�_�,
R�D���eB�d�4`|��TD�vk��G_���(N���+:@t���ȴ�Kù�v�U��<X��χNB���t���5�,H��^u��t8E�%�Y�D�I���
��ȡ<y4^���"k�
U'C�Q�x�������-�sA�J�s� p�|I�p*~��P����If����݀TtK���੆���;����;��-��w��CG��ݹ�����G�]���IX
f!��0bU���I�C��׽o�I{l������8|�tռ"e�5H�	���^8G��p���c%"��*gt��p�+�SAs��ȟ~A�P����l�xH�A	���y��`ǚ����y`����͇6%�d��X�� ���-�U�e'��A�H��/V镊�!��¯��Ё��U�^�t��S���x=��(�#��_o#U�����:�x?Y�5���ź�Oc_���5w����XՈ���$�S�J�
�E�UA_>d�
j�%M;�ʠi�zF���)����(M�d��)�㴓Wt̪`��)#���m�g=����(Z�}�K_vXlxVHYEB    3d43    1030�g���Ug�bZ��O�5tp�bF8@r/Ҟ��pߊ�:~���n��͢w����;+�d����������p=�o��<�v���}U5�X����ܶ_;���i�����vեL�\�/Ïbw�������� k][W����/�ޏ��Ec��W�R�T������@+�Q 5(��~F���B�υ�a$e"`؜%��z`���?1b�Z��P?F�i����>��{cIҜ�!�;���kg�֝��p"j�G#��&���:7�t-й��*�����mf~ۀ��n��B�t��롑G����~�a�J��N�#����$H_�I�	"K�S��_q�'N7,���MW^hq4Qݲ�(ց[��)7)g'�Ï�\��*6܉�ɻ��<�S��g�c��{ ec���`�ı�C;t�i/	֖�k7ݤ�U5��UGP�[͊�E,��,Y���ii�Z��+l��;-���>ꆙrJ�@Sn՛u�[.�E��yE���7�}��v���(�'hS+u��\�A�����/�VwП{��x��!HTa���uA�K_��?Q���zR�����_��x*Qh�釹��B�������ls_�T���/��X�&�(��-��W�����m�z�j�J3�Q�w(��"<��3 �w-v��S��Fu2�|�z-��?��HD2k+,f�z�\Yk�u��z ��g�6_�+�$�J�Hb6���k��	Դ�!�˸� <%�0=�����밝�4�J$R2�1�
�HGI���@ٶ� �
x���G<v�qo{�����L��`�,F4!��չ��-�*�cX��p������M@׳bE�Q��e'M�c5�\��4�k~�d�0��o~/P��V���R�gy�S�]�[�T�!�W���3����U0��1��1<0D�A�Ĭws��_��O&�:!
ނ/�t�X���9�ޝ���C�'�8�7AP��A��D®hfנx��3���0�v귦�+�blcД���abW��l1��r�<�7V��|��J��S����eMh���ح��vs�i�o���j���+7���=�6�z8��F�~l2d�H�ޚ
�[�,ꝱ[j`����7���qա�/Hf��A���5�0.#W��t�:�(��X@m�nl�����0%|��sCo �z��gpJ��uP=-h�#�a�t����� ����5��8����<Z	�И̠3�笵��⚍Q�Z��������υ^�:1h�b˃�R�PT����V Q���h���f҈��SR�܈`�)�m�w��W��9���娧�1,N*R��e��j���%�%d�{�Y���/YqZ,}�� 2s�Zĩ_d ���#*cn^���
#&�S@4t�pi�\	���w�@	/��Q���+��Nl��(����0��ge�����Ц�Sۀ����V�_ʭ�� ��r)����I�?��)x�޸ܶw�:�Z,݅I�$��ŕ�H��������1�6�/cG>��!��Öh�E�"WY� ǪQ���i��5ý0
���8���ړ��(�Љm�G�v&D��ֆ��Nv���J&-p��"��z!aϑt���9"$�uţ�д\m�R�ocQ�e�x�B�3����<d����*���ڪ�	���:�D��}��;"���?�����E�)ې\�2�Oǯ0�{vɀ0�}0�n���L�@Eg##�<F����3~���֩�<Q� q6����\2�X�Q�BnmcU�&�NQ4k5'�&�ϸ2�Fx`):��#�^痃"(�{$}��XD2��#Y���%��׿���;�fz�Ը������@��&uL�rH�D�o$�'�'��wTΖT�s(h���m{q>?�?�HǞ�������K����i:��U7+J�H���D�R��<�j���QCCۄ��ԗam<k��T�V1�b
�l	H<��/�-���f��b���&����96=�Mc5��9�#�wJ<����KE����(�@�(���}���D��	�#@xy��n�W*=��2�Xm%1y�G*�# �gui��j��e썇5vle�ʈl꤫R�`7��^��\�H����lsg���b����#����U�7�Bu_��d�n:�Th/��
��H�����+,f���)��-�z"��)�Fͺ�`���5O�����n�ex�a�(M.�c#�V��{��#�mJV�BRjjA��p�@��T�zmG�bc�.�ښ��~W%�-3&�mml�F�6�
�.Sۉo 00�������[>~�\��"g;��.�(X����<��잢��b`7�g��|r֊�A��c�1���:0��Ϣ���J����wR�M@�N�A"��r'���V����G�Õ{���M�濺M�_9�Q�؟����zzz���`F~�����Ӯ?� ��j�[���b�0P�]E9,rl��j�e��f��C6��6%�6f�l���̩6fT�0�iJ�`���mg�8�p������R��!Mdo��jɰ��?bfa%���:���ذݲD� 5w�~vL��-�'��h�W%��t�S.A/�1c�p~x^��a!$�#��qP<\<f�P4� q��v%�K���en\�$� 3��X�C$���=�I�i� �2j���Ĉ�R@�%<訳Q���9�� ��h��n���k��604�Ϳ3f��\�=��U��fyҨ~ӊj�c7d�qD1fy���N-�㛆c"�iQ���)�m\7c��\9���>'䒣���Z�dmL�$e,�m-I�4WI��(�7�B\�a{����9����=��tJ��1a��O��&�XS��{|�Q4.w��;1���bCx�q�ڵ�=���G�����pf���@�Zi��;��M��ho�����0آV�k�NǏ��6�3�c�3�4��w4x�Y�ŤIp�Ow��@���e�X��
��)�4K`�f���q��3D�me8�v
Z3s�.�t�K{�y�@�Z,*���h��*kx�]�V���yUƧ��6v�0u�L�K�}b�.^�����:���.&�,߿���dr�^�	$�@��PSX�0AK�\@Y�}o  ���w�6p��NN�,��A*�f�t�lp��7");�y�PX���j@�M��5W�*ٕl�ȪD���mKc��V�~�|�h�J#�z�?�Q�0�'�Z_w��t��`��|x6�-@��h��Ҷ�]����zJe�Ő��WL��1��q�]hu'~&
H#�����?5G���С�T,jN���P�>]<�}���l�D+���'��߬�Z��6��u��dR֭�7��T�h��G%�E58
��L�ZZ�\�V���^�:�&q��BbK�����5��K{=��eݶ�H��P�#9#D|�غ���g�i-���
	�X�Z˷+�@�f��Z  -�_���&��:���:"�����6�B��a�N����9	�x�����w������4��ɔk4Ǥ�̿�[�`_�hv��z&��&L9�!�-��(�L�uW� 8���4}�-z n>���S�,�v���$�A�qXؾ�D�&x�Ef���v�B��ݨ��Ljq&B'}���~9�n~,n;���*�R��b-&����D�� �Q|�}ט���Z?]�wӷǖ�*�;����&2(G@���&�B�j����~,��\/$�G?o��2����
�4��@���-��6���џ.G�Z�p���	P�v?({=��~���A�Ռ8 e��Zdbլ92�(1Ђ�V�1ǡHŽ���������	eT�Z�.|�1b�V��º���Z�t���:�_��=�|}�Cȹ�({�,G�Ũ��t�-�)��B������%�nbp4x?'mFwf]T".��2�h?mx]�R�[��B
!:.,<&��")���:�6�'?��wR�b��
sonNI�F.`�F���E4g��iŉ.�y:�4c���).��W��Z&�%s���5��nb�ܵa����Ӷk��*T����5�1������4�j� ��5K��M����oѮU