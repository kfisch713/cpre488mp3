XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���'���Gh�=lpZ�����R�<���@�R�ۿ���Y�FH�'�=�����"�(.|��4��h2L�[�΄�^������:Ef�b �k/1�А���:#?OH�_:e �.����[wHj�R�_夸4�lO�S6؝�����Zz^M��cў���M�/$,�;��<qf��{l���n���O`g��3s�l*�U�Dγ�T��>��9��챛lF��ݒC�x�����/�O�W N�����(G?Q��(�T���(�RJ�H",�դ��m*���ɟֺ\;��N��]Q2z�r�'� "Y��&n-_�i�yE���oF��V�'1��=�Ħ~��K
������%%$n��1��+�� V����o7'��dA��H���C�ȕ�#D��f���s4Xq�䱗q��~@�!(��F����@�q��\*Я:�����7��.Lz�����:�\Gj|����٫�D,2>���dE����c��~��N�LD��Z�os�ى�D�GS,O���S��x���a��@�⚩8�pr�/|��}�w�B��XV!+�g:�zY�i���i$TH��
�wgL����!Z��T0��CVɸzԣ�Fȶ���N	|ۆ��nԃ����r���j��L�/��q��+��L�^��#0��c��%�ep�xhlZrM��+g��	?J��!d	b8�M�K�І+y�'�O�?H�bM�<�`�B8&{�ݭ�(�'�L3s���wAlT��R�oOOeW�[&�{XlxVHYEB    2326     980�~����nY��!~�F���@F�������a�c<��8L��:+���Jc�H��Q�/�@��)��XaU*��{��&$�S����=ò���K��C�|��
�.�3���Ϲ�k(~�׿<z�e�p�j�*z�ʫ:%��EoV�X\�=/�������>
p'��ܠ�yBJ���OQ��a߇��Cqy�yh� cf�֢�t"Gxg�}�t�8g��1���m}>�
Uj�Oqʄ.͜��L@�l���X����^;��@UO�ю�U-��LD^��9��锱�e�'�2�4�P2���'�ُ3#���]�^mx�.>1O����"|lu%@�49W���J-�<��<�k��~D��	*N�G�g�2��C'�z���1^p���h�Z����dP�;B`t�G��Ƿ�y��u�O�JcLI,E�(9���I{�;��\ƍ��
s
���tˋ�L)�� .��q��D���
u�}���ʏ�2��֑��^s�0��Ι�+C��}n����I�V��k��Q5Hʑ��Ɉ.�;�� @%^EH�;�ځ�^n����Ҷ'���
��pG$P��+�����]P�
�ޙBN�w�afI�|����r��=M"�|k�	����xu�c-N��kZF�9"���^��p��z��lMx���x�(n�K-P�%��n����y�G�T2U�����8�����M8h�e$Um�`��	��������ʷ��4;�D�!����b���h��{�,��i+:��J��!��}[�S��X���7o��C���@߼�Zt\�}���}�`�H�N�h�^43��EAҚ���&ɏ6�ye��}y}(f�y���f(�g�89>	�[?W� ��¬֕�	1�r#�(8A����x䱭�$-y��ľ��J��dВy�=+�\��AP����,R��<�=������h�y�ڴ�Mz����@��Y�UJ�{����qai��M/�{��^]ȕӹ��GĮބ�w�՜�[d/��7R��P���s�58U�-C���������b��4�}�����X�Ȁ��y�3���6�h'm���h�E��p'�ANC=˜[�bكE�H��9I�8|�|a�A9� h(�׾>q���o��Z(k#�X;�h�d�؁m_Mc^#"��IW�RG���t������u��.����W�6,'���
�m�#�H�(�w�����n����_^�3����i�V�_*�)Ӎ��$�� �m�/���빡��1���i�;Mc����s1�ᮓ3�'�֏�í1���$��5���YRd�M�ؘ-\�����Z����	|�򾮭�a�MoO� �����4�����'�r��S��0�X��:���6,ی��o����S�Q���p�t�A9�aJz~f���/�}-vD3^�ŒD6��+�58�L*v*��~&��8%͓�B7���B���R����!e"-�y��3���{a�"�|�����
ӝsŭL�ֳ�wC'	�}��MU��>��K;����%wL��!���df+�Tܥ�z�آ�SV��a Q?p[���L!�������uƣ8K�O��`�˰C٦�g� �,TT��Хa����o�q�>���M� �X��?k�"]d8mۜk���D19������w)�sH�4�O�9q�&�0��D�y��{�m���"��}��Tf�'p6����F�������<�	�����R=/�,�9�e<�
�/��!#���wK����>��{���<p�/�1�=Fֹo�,�0-�K�0*�vr4:�;	i�l���U�4���ip �E``
�7�ج���D���g�<-��? $�����S�Ⱦ�J�5]��{H�ٻ�8�B��DS���˸�PL,<��⊮Wqp��GN�E�@�}�Y�>��2��X�X�p3y-ߊER"��Gu��CY�.,��C�e\?8`u��O,^�,~K7��X@?�4���s�����~����f�w�L���O���rN����Ӫa�=s��P�H��;I�X`I-Z7�|�k�ya~i�B鶭+(��~�-n��Qu��F;`V�l��[M�ZnvoW��_�l&t��|�L��t/۲�:Jos۹��9}�	AEŭ��Zj1�u���~Z�i�c�j���6�͜��S8�
�����V�>��|�˛MD��}<FZ���̓Jq� K�@�ua�e��-^���ڜ�OI
�1��E�b�O����5c�L�9C�q�L�@�O8�G�Y(�͒�: <�W���W�W9�qe�\��4�m��?<#�a����8	�H�f�^��+��9A���	�̸��vLv�r��3D=�DX�;����������m�����ᣏ��!���	m�7|��jĺ;p�tm�"�L{0�U\���