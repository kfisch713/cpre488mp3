XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��V��
��ō,z�����J���/��)$�m�A�L���+86�$|�7t�9�%'��w	�o�
g�$M�8��%�^�ٽF]�=D��
<P��e��O�}NԼ�	Ú_D����B�c����%}���^K3���Z-��>f��CI "+0�t�p,����6!�BŒܗ퀠��i�ԣ�[7��`���Lq7/�2����;�	�Pe����"��|�-X��8TǾ�NPL@��,҆���;m2<>{F�\�;E�����H(P��7X9d�'/)t��,�� ��O$߁]u����M;�+���Ϊ$�d+�G���ݹ��+��U��߬�x3@JW�f��pф��t J+Y�Z�s,6*pÆ7�����l�{���iu��b/���M�go;�!Є� � W��}��f9"j ���"�J���C�{�n���_}�$��yos��&[��-'Uw� �2�1��ߏN���d�]D'��>s����Iǒ⫭�s;�E3������P�mQ��]��:�����O�ٕ(�ߎ�oZ;����p�3�و5,Sw��Ǭ��U�^�X��ޯR �MvM=@)q�yi�ƺ��j���i�-���>{�}k��I^�W�Pp�0l��&�hS�yt粬n��<����?�9Z����b��=ع�{q�@�˱� .�U�'����#��缾�l���ʨ�<��
AM6�{������ѽ8�N�"���DV�y-�B���dR=�b��`r@�z*�D���ق��3�7XlxVHYEB    3da6     fb0���i���ϖ����C�[���@f>��A��Ą����M&�U�*G�!O�~�B� ����s'qI�C����>/ò9�:�4S�&��Ͱ�htC^�P����*���,Fn�X�q��&��N)bg���Ez$�Kϵg$���p�@4r�DA0aN?�\�$�����]�7���L�}v��ț>���ega~�`8����?��������A���ځ��6�!>-L��H�x��;�;�s�u+L���S{X�,~�	I�l�#~�TF0[��ev��/ֻ�'BM�=ђyU�����m�XL��P)����6���J�T��Г��F�1Mǌժ��;���P�}ES�;�C��%���W�M$���+�\*����+ZV��)8\�B��u�G��Q9N�ؚ �)Nb����PKe2��xӘe}L��]k���q�2/��썾��|���H��$+��&݁)!�塞��u�.z��_M�6��,�ĽQ.[~�s,yf���T
�\�"7���rT�㖴�
�|�����c�8^����p2`4����*�Z��-iEϛ�;���'J H�B�`1�ӵ����6�7�C|����8�]]����&�@�v���P���?�H(��{aeT����T:#R�����F�6�*���� ��q�?��� �c�o^��a��f�@��z��%m%Ye����z�W�[�7��l���93X^5tV3����[!=&:U�V��[嶒;ɸ}6���J�x87f$ӱ��=���DH�QQ�Y_N��fVQ;�y�������,��3kƼ��Bʱ~Cx��S�~.�#�|9'"5����8�Z�I�b��Y�P�do������V���%��d"I�7�2s�V�j��GI�4��4ǅj�1݂E
�l��r���mַ�' �v�/e�Ci�vW�9�67?��=?��t˾!N�>?O��{����^I)�!=�-!%w�Y?K�PS�,��f>d�5��vӂ3���d>�!���`�4t�����vM�����-�H���������9CT0n�l��
�)��
�p�!7�V}j-���Q͡*�t�@�BCD�S4�b$v���,#(\���(�2R2]�r�����~S��!�_��J�c�xA3(V������Dg>�|�]�@���H*Vv�l���uO����D�C� ���MWK�&s{J{����$o�A5�	��&^��J^�R��lcQZ
�5A��e���V)1��:3l����Sw��x��X�Z�Z��Br���-��|x�ܘx�:+�G����j�l=~��M�J�YDh'I�1�g����-�5��K�����7�`�B�������U���p �\�6t�"�ˣ6���ns�����^ċpՖh��:	��&�1u�ޙ�������+����&�bއ�òh���M?
�� f#)-Z�:ˑ�\2�Sc��ME��h��v�0�K��P�>��z��"��g-������Zw2ӆ������1��$I�z^�Xn�����nm�5DE�#܌����xn��%��&���x�u��Clg�=�[�?<!�d��H���-��7Z�,��/�HO�bp�޳ �����`~W��y���B^�q�$p������w��^j]��7uD"׬��� Z�t߰��=+~r�=�@�s��3ꆲ���J��c@���Y�6�(��a3v�wبvm�����_.h��ln��K��2���!!Z�{r]���KҀ��O��P3�"E�J����D������)�P�v�Z�d%��8��d<��N��0���L���:ێ�E��-�:o��ʁ:�š��כNw ��D	�n���f��^�A�eg̀⵰�N�(<�� #>T�i.���ArY
��Xu���>��ځ���#���B�7��e6�Ťf(m�������ڄ��zV�$}+�����;�Ҏ*P����%?�Lhq�e@5ړ"�h��\8f+t&��]L8+'B'Wy���z���nZ�d���Ӓv��)��s���+h�6ݳ����Q�B�8j�%#��XNO��2SR���o�O�C>B�б���ɾ[y,�an�/l?��O��. -09�����(�|J6&��9X1ʼt�{�3B�8������9�n�E�Or��{�8���x�C2��o���G�!�?�6�c��)�wEHs�&�q���{d�Q�M��	��܇w�\(8����|�6��7�@!لK���0(�-�E��g'ɞB�iۚ�o�/O�%t���b��U ӑ�9A0������ڃ(���PP�ؗO2����d���,�=�y�I%��SOW����P3H���� ;�g6�ƅ�����p�Lg��k
�!/�H��H��C{[A|"z�����*�6/����K��=�U=��)�����MI`����y��g��w�^�d�S Ho��Q7g$��&�P�2V�B
nh� �=AY|,�f6J��ơ_�R�/��jl��:P�ۼ;����]Xv�EtU��e~��RDf�����.�Z�V�8�ڙ8|��v���jw|�GR,�iT
��2��N���$2��މ
���N+�ވ�"��0ꟹ���V�_G��u��!|�F�<1N�Nf����}4�p\��}F�A��bC��>qו/pf7u�V�J:r�a���wҭ;���G*C.�FI�q�"�+�N]�x���>hh�Q뤜��*@hl������J0K9D�s
��K���|J����e�#�p4��3��4!k���ƛ�4z�3��Ȗ�zXB��cp����v>rJ�c��|���,c��u��\�4������V�~���JשD�j��E=��2��}a�yz��9�^�}b+�aP\oC�9���WK�s�� <�������&�+Y �ƣ�Y��0%4x��2ً6��,ZS���I?O�m�MW`~b�8�p��C�e��K�w,�byH�w���-������)w��T��8"f��kD��`�(?o��z��A�~�Zf�	۱��aX�h�f���֫�B��/'X��`1�߻\��>|�"��w�Z^4h���t'�ND�8��;���L�v� ybw��T�����w����j�*�O;��æ(ڀ*�b{mf,ք,Ϗ��%@�o�z�4��c�5��Fq�������1A&G���G8�3���͝�bɭ�)e�_r����؄=��\���7b���� �T������W���hO���<BxtKVKE筍��N��Z�����\�eJc�-C`avI2��<%ֆf�'�ie�]��骞@����F>�A�P/����ö+��k��[�;�s��s'���4F�}�9�ć��w�[[�B���z�9��=Mď�\�N󷥎�ٹL����4g2�g���3,fk�Ҩ�>*���,�_�G��_7P�=����Fhy�hBR�����6*�3n��Ȁ�AÇ���(�I��"5��&5��#�/3KjW�9Yx���\����\君�'�b�����˺�� �m�DV��	1���T�f���_���L	��&�L
��q6�`a�rb�?����Q�	�gb:��cuRI:ܭ�C�<���i�q�D��
M����. ^��>��r� �����_�q.��=H�'2��G�'D���$��EeL�i�����@�y�Si�|�N�x�����=�'4��k���/L��Ҿk��u�J�&u
W�5 ��0Z�x��X���ڐ�1�H$!�unC���N�����a5m$�aO�:���l��ܲ�B}53�����%S���H<o�����g��A<��� �+�*5����i3�o���Z��T<�u,r�/�����c�����!w�zC�OE�8��Ѥ��VVF�l�ޠ�[�L��