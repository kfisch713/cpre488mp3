XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��8�钆�J������q��P�r1^��7'�J-��9Gݦ��{����h"�ٸnUT#̸�c�li+ rZ�c�ȑ���c}ez�l
RM\�x6�ב����l���t�v>z��о�Nt���ìt��:���" $C��ņN��.��sm�څ����Irr�૷.�z��"�S�w��ٶ�G�������bo^�����m��4T�$�9�	WKq���*�%Y��w��+�i�Q6�{���m�����I���+����XRؿ`(��ʉ �c3?<&D��S�b!>cƻ��>KBe�7|<��kÐ��7���j?;�Zt�O��~�I���Eا �������>�ˮ�TMC����P�>�0C6"ȷ��eɀ�3!��x:��CGj����Đ�f��ͳ˨�]I�\OOR�>�V��g�C$O1XlTS� $��K)�/�$���s��"%��t����o4X(����B���H7V��2�A ��(2m-�{���S�<'��r[~�B�}̈́Ǹuڴ�D�k�w�O9�����3��:�?x�AN�m������5��О�p��$�K�5̊k�j�,�.ťa/A[�l�����<3�2oo��:�+���)a]�a����i��v�*� Q�)S�ͥ�#��ġ@i9v��s�)"[XF;~~d�K��ձT4�}^�)f��PX��pIaP�2���6��"����`��||W3���}W��d��)��WH�iCr��<��ʥ�FXlxVHYEB    70a6     b90��U\bW�DO��Mc�ѽ�S�f��m�--=�i���1�.��?��Uc��27�^�i'��s��9��ס�<�BGq-����]��,Lф�*ފS�%�q�#(%G��bM��*�#_{��I�C��vF�c:�����0�C}�������N��Nh��p�_����:If�#��ĸ�����j�2��3�6+�Z�h��]���ˢ'����4jzH����|��f&El:_�q�	�s��5x�ɤ��v����J_p-���w�]�� ՗�Sv��1�2���5?�N*������(��nV�Z�!]�"��.s��p/X<���? �9^�-����̏ol�gUk�f�J�W�l�q1�g1VYp�V'�W��`�J����q%��~�ZI_ũm*Ƞ�MMJߘ1�
��!���qY�������R�Gl�C:u_>�D]�vE�M����Z fSD�V&�k����4Q�˾������<1q1�d�SO	�$���qa�(@QDW�/F�۬����f�-+F���k��~�jPSP	Z�دl>������;�b�b��^W�D����Q�b㔾A�����i�9��҇IR[a�D$�%�����_�t�}ЪVkzi��mw��A�����D!7	-t:-Eؚ[w����iMd2H����0���� �y5ݥBmԔ0q>3��ޜ�����x�̢�:U�!�-�f�9#R[��U�[iO�>U�,[��id2���{�<M��GO��bA�qe��Ċf�6 Q�Ԯ?�AN��K�.��տfR(����]9��b��D䃲���J>��Q Y�1�̒��)�u�!BU�}�R0f�}?���dS��;�	�#W���8L���6�5�ic����d�����������i�6$xˉ�S\C���L]�38T����n�Z�]ad �%���H)���X6}-,����VK�Z��nLo)�������s��B��'XծKL��a�<r�\����&��b��3l?l�sPm��Q`���H�ez�I$�}9��p�E* Q-��6ߠھ���bb����@��i���19@U
ق b�Q�Ӏ��ۈS��k!H?�c��^t�iV�dkx ����D~�(����y�c� ���U�w�cYw�����e/��S?bcg*��^��8k�{M�~U��1�9���x�T�|;?�K�e���|R��|��\��φI���Y��G*����N!�����'?nJx_~��z�z7X��a��u�5�]-�s��kʄU!h����.s��N�|�1Q2TQ�^��<7b���0�
'C����=ĉ�"�@���x�I�A},J�w�[lO��L�윹9%E?�ҤDd-��ݬ��P�^���R�D\z]u���u�n��3=B�VC�����NW��M�Ռ�����f�"]}�2� �Iep���&dR.�$�=3�w�UT������k��7�,�aЮ0��[�H68_���m�.�9a�9,��&��e/ҤC�Ƨμ�F�D���ҋ'�9F��\˻�4~���ĖT 4�e?;G^� Y�G2�8	l\`��mF)]�k掑Е�x[���sޓ�+^%��\�`z�^�������}jS(����-
��N�p��(h�!�����X�K��S��g�Z6��7S�(x��T��V,�`uLD��6�=atrƦt�0��E�D��K�:J��gWef
;��7�xW�WD$��)D�ÿ�O�l���:<*�����텤F(;��EG�F�>t�
�I={+�����A*��d��]�7�mSwR�� u왶� �@��^�p!p;�?����＠*�l<ذ���UO-�`XcoȘ����U�wxc����B"��� ��UC���|0B�%On}�Y��p��Lp����r�C�T��[�>�*3Wz-[n�S��Oe^���g��6ᶘ'��m�/-o�'X�O"��֚���*"��W�Fh����~��D�(�T��I�%I�
��g�9mc�B_��ثd����4v�s���JI6\�#r�U��[��?O��
��D�\�@ڭ��`���M�7���C�S��{�2�5A�YE�#�M� ���[&g�=p��>�
y��;SC<т�Kx~��5�}pJ\������\���`������WM~��ag^<�t˩��بu�zŵ]�KԹec��m��duX��������ч/�`�`��Pβz>3�ۊ���%�كs�XxLj�H�nz��p�g��#ph����;b �d��:��}X)�)�}+��'p}�h[C���Pj�*P�L����F���X��vT�d��NQ�*�x24W<gw ����Ũ�uϑ�>9#6�&Vk��|�yZ�r�|e&�� ����x�.�������rB9�R�z,��8���ױ(7������Y�,�:�Ҿ��Dǐy]1񒬴1Ӛ��,c�����:�ct2L��3�[��$��qY��DKe��P��I��T���r59wK��)�I
��Qe��IE����ї0zE冔`m�U~3̅��t���dэy����jӦ�\�~��cI���V�H�*�r�}��@�m�'[�U�%_�}�Ө��J	A@�@[��H�!�����m�~tNZ�<k�tY)����9i� o'EM��1Tc/QҦ�LJ�x��J�\����	��-�4�kʚt���'׉��XW�9�YU�Z�{3r+��	>Z5������d��p�|Ꟙ�v־O[��v��"\���#�����乱����)�vQ�Ɩ��O���+�zw�?����i�x6�a�ː��7f�����h=d[�y2�8CB���?���Ԣ�A��e�v�Ʋ�m|e���hz�U&p�*T}�=�{=W&MI��q7�8��]_L9���=