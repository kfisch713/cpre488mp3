XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���Nv�F�Od]s�ۂo��Ӣ�F�?��8�����ob�d] |i�	�)�Y#���n^�`�t��t2����Qv:�s>�+�/��`uX�H$J�;�ݦ�'�v�F�u��yI>��p�F"��۔b�8�b�R�>�ѥvU�-����W�o9�Gp��3�Y�I'��7�Zq�!"�ԧ�������wT���J}y�.�$=������X6��f�i'���Pc-�]��'����=>�$`��}��c�z�]f4B[-�쌆�>��G��l]?�f�Oy�V��L$�$s���'l�t�F�{!Ǹ��I��n֋�m���nD_R�yM��>(j��)���sj���˘w��|������]������ӎw㈀�p�Vrf��~-gIw�a���(�̎�1�g��3L�>�Rf�8��$7+���O,��B8��f���Og �@P��v.�ޯ�@�:}8O%ק�i�4^��O���'�v���Mb��A��q����\���ϻ�[XR���O�����;E@���w	�.Ο/\��o���_�-�~�����2G�v�|��J(Qa5��.~��|����N|
�ӗ��Z��pEAY���Ml�41�^8E^����婄m��GVMl���7%��qR��m�c�����B�},gN�'�'��ܸ��R�)U��T_n�Qו�+}_��ô'�3R�E��3On��K�zb��W����(o�wue���M;*��]�F�O���D��X�`���yXlxVHYEB    b087    25407�����r��j��Z���3��D�j�%{�&���h%����!9
 ��vX	�@1	vS����Z�^n+?�4��/�D��Ӟ�`Z��z ���}���l+'N�xi���7̨�ZPU��3�j܂$�Z�Em �#�2�Q/���fԇ���5q��HZ��|lV���S�K��޻.�j�S�����(�Aeޫ-����څ7W�awO0��k���L}���o-ou��@����tKlj�{"�Q�����	l���ʎ�2���C+d�g�e_j�&"�9�$�����k��|�Q��0~I�ļ�J݄�l�J��=�>�Nj�5�m�\���fKJ�#db�ϛ�&Ece[�k�D`Ҵ�ݛ@g��1�D�d�"��9� x�!g���T��/�>e�U�%�.�`� A���P=��Շ����u�=��*�/*�n�Sf�����#�����]�2��QG�;Ĩ��X�{k �0}焕��-���tF@o�Ok�q�w�ԸA�&(V����3���T�F�/{=����[��[U|�j��1�W;��~tQCH��
���4}XS�N�<�8�f9�^S�����j�,��riR��w� ��)��$C���SyN�g�2�����ɝ�j�>���\��&�*���^��?3�"NL�n���L�vI��T���MZ�I@t�g�i_�P��	�|�d`��<�G�؆L�JP���R�p<��+����/3"xp� ��CA��?ǲ�*�5�{h-��iq[�Dr�H�A�W&Q�e Ԁ��u�!��!�SjBܵ�b\s�����&W�'���}js�59,F��Xw����#A�+��ɖ�f(�y�Ef�'�lOD��5���2y!	l����<�[*N��Q�80�Y��k��,s�y5>/w)J"�s�(���Ouޤ�w�۴:.���V�Zz��u��S�-M\��|�^�DwdA�b�B�IA���"w����];.|�Ě���-7�� =�B�y(�ٲ�k�\vm^�ߎ��18k��4X&���y�������=H��C	{O����f�ՠ_J	�%@�Mq|`fs��&WAĨ�$��d_�ݐ����D��6a-���#��]D>�������&#j�	Z�fn!<����퉡��Tn)�z��wq#��1��}Z#*bx�}����%�Vb�hd[�H���4��ӗ���|�r��/SS#U�2*\J�����T��-	Q�M�\|�����n�xp��/�$��=�M
���2߸��R"`�q	dU��X�W��1�*�*:|G +���v5�q�GB0j!,?v˟<����{Z�?��r˲9Ş�G�&��X������C�NE�lW�G�R�y8���L"s�x2�U��ŵ@@���Q���~�+��}f0�LUS�k.]��O�b�nB�b�O�+�~�������";͍�l�*]���VD21ض#�>�����B}�Q-���������c���QX����1\����� �]�T�]v�Mqv�����wPaL|;g~��/J��U/��}�D��-Φ�ׂ�K"1ɠ��-�Ix0�q�:��o᧱��p���a�ߣq��\�:����4��&R�E��濠�H�c��%�vo|�q0�����Ӄ�<�<Ϡ�77=����bF�g����v�kG�f��vX��(��A�_BBjqp��S3H z��??�`,�"�
�?�Ē��g�d#qƿDF#�%�酪g'�=�X4		��ph��G ��g�����,��{C����
V���NB���>V[8}�'��Dlu��l��j�`�ƞ��<
ҍ�y;�Qw9���į�I4d�U����?u�Q\�MT�R�5)*�Ʀ��>f��2�6Y�E��|�@^�~`\l|�a���D����:�J^��)�de+�/A%�S͋�"��vټ.G�����xvO���	����m:�7|<����@���&�I���/O0��o��Z?W�9�s����%Ye	�_oA�C�w�����HG�E\.<���A�M'Q��=��δ	(w����6��y�I("UVӼ�͢�G��a�h�f^pJ��Ğ��c��Y���K}����N���]��;�ݪ.%��[��i\��0ʚOc2��h6��k��"<����uk�X�Cv8?
�j2��Ԏ�=�;#k<Cc��v!� PH_�rMH�țx���	�x�B���	D;Q��n(�d��X������a�q��!��L���t�8C�	�>�(�;��p�;32)Dm=�z�H�*�3�
	��P��=���~n�B
��t�|�p�0F�4Oڇ3m�τi�k~q�.��棗GT�83mw4v�7�8yI})�0��{�+~w�7j�I�'�+KaŚIS�lG�^�Dj�؃)�)L�ה�`*�d���>�1��_K,Љ�(̍�)yL���(�p�ւ%p�<G��\5|77�{��a�@�w���,���Y*�+�Hµ�2�������<�J�?1_���M�hJwt5S�����C����}����	��&��{�u���E���U�yK�iʆ��+�
�ɫoa�_��o�^Ժ�X�g���΀6�E�hy'ki�;u}((�a��t�`�9FI�|���?�QT���W�
~���;��Hw`k?��D]��i8`-n�vվ7����#�Rk�@Y3����wU�0��/J����A~V�nX	�+b�XL=3��ga�I��2A�h?3�Wۻpث(i��!�0�����ӷǜ4t��C�i�$@�=��O�4_��W�G��Z�q��Oo�lY{�ELʹ�V8�	��c�뗤�Yl�Ou������I�8s��}�2쒘��]�2�\Dg�TG��Z�"shK�W�.Q�@,�x͹#\�HL�|]:�si�H��W�{9����o�1���n��_S�=�|Pz���֩���M�-1�M��#���J��Xqx�Ɠ����t��l����p�F���[i���~>��Y��4��;��D���>/R.���W��a���x�!��D�]�!:�g��zYM������ӊ�|�(�h���l�~X����!�m�@,�2����n'V��Y=��ZK���H�n�i�l�wl-�Ve�2!Ƭ�W��=���Plp��� j�Ry�4�V�V__0�nXCL?�;k�

Fa���R�gJ�eK�������m6��|[q�c8PWM�(KQ�h���{w�������p����^�`Fv�(D)��۹�>%�e�E��/�?b��k��}'�OV)�����z���bw���+6!�����db{[V�$X���n��,�&<?Z�n��/�%CHU��i���Kd�0���k�m�Y�+A�$n�m��3V�a�
P7�B40I��n�� ��h�i<�:0g��敍�d�NGЄQ���:�A���7�es���ɥ0���#�	d�i�����PG�����<F�#��"�t�9��zH>����ø���k����(2��2t�\M���o�[8��:tt�����{��(���p����W#���3}�d�$�lh� ��խv�?i4�f�,���b7r��AC��b �}%P]�vW��ʉ��C;�ف�ݠ�T��HT��י�~[b�e���b	Е[��7Kݙx:�r�9�P�[�d
/�/��a���Vnr�A��:�����,`���,`��*�7��Y75�����-��Hh���"�_W�tJ~<Τ�D����F�!�F��ck0'BKThx15��3k��RS��X�5�Hh-��^J�M ؐ\��cR��-�L�p��{�����!Y+ȸu� A��p���EP7y��Ai�`���t!��������b�
�-�f���� b!�v˟n��,�+y�lSm��c�ҫ�Wwx�e&�OФ�&�77ڞ����zf�)��>�(�B6׌�<�M�\ H1�ۺ] !�je0�TuN�Cx�����{m2�Թ�ӈ��Y�A�p�sI&��0]6y��C>���+�5����\tԉ�(�K�ʼ ���<���}���T �8]��ٟ_��� _~�TDz��1���S��N�'�Uk@�(V͇��yo&K������&S�h��ffqN�vQk4!hc

��sI�<<�.�vٚ4*�U�Xf���uy���}k?�[S�EJ{���8���Z#��,�E:�saM���>�Fw'��������ʍlyŀ�~��w��#��g�8����S��困���q~�ޫzX+�y�-�J��k_,� ��38�׀��� �֊��'f�F��P���k5¹"<' ��W�D��>5�z�U���B<�߸Ƿ����7��q�p}�Q�0E�?ةh�\n"	%j�R�Y�K���C��?`l��\Bl��E0�����a
=��6���������*9T��O��RZ�ys�Цfw����S�|p�(4!��Ue��ʖ4���<�@cc���➜Ј�SËĨS�k��,գ��&�.��ݣ=ᄀ��U;`�6�������{���Ewý긛E�_z��{Mpӧ"��j���!S>�K=Q�Zn�Q���̜��)�$o�"KF9�6T]��*']�P��Aǒ��p?�4Ps� !~6���t�V�ϹT�$�"}���u��K6��3���x��H������FV[�Z��Ǌ¡�;x
�
^Ú�әR��d�[�Z����8D�ڸY��`�MmY��7�7'�+\��'������:`߫���Y>l�?�>!U籠��u�h�`Ƃ5譪�K��)���(:�"�0�Pd���J<_"!�ň��a�t��=�s�t�����@n�D �7��~���-�'���$����Hv)���������!yE�>��O��:TlƧګ����(Xr��\�Ԟ�d��=1O����|mxm䋸\M���4A|�	�����;��|W����M�9/�p�n����Ȍ0��۫�B�=cg�+\-*�CO
l��%��`�)���5�9������\�Ӆ�9��L-_T +�I��bP},�������1�$�E��;o���H��y4$ɺ��6�E9��0���l�%@�B�dU�M��E%�g��h�3�ʽzX�d%>�sZ ��%s�>h��A K�'�D���@C5'71.=�#P\��c��,p��]�!���_8J��:��::+dL?���U��"���b!��ì�y�o6��A��j�����V����+.����Hs�o���}�F�t��,�t�_�S�sh�Lw�{q�P� �C�*5��8��.�]&�!��X��q�Fj��s��׽�]ei���Ciy�CX�>���b��ޥ����Ns�'a��k�ɜ��t*�1A8L�_�Ia��RQH��xVBFevq1|g>h�0��}>����ة�b�gǩ�ll��@ЯDY6[�F}����i^��q�2�-}����s���l;ms.��Mm?�y�`'�ϖL�a�����8�5����+�2�O��u��Э�P5V�ij�����̳�<�o�fm%f��u3.��8g�M���f<Ô�o�+����\�ml,x��WY� ���*l�K�^_uA�P���[M+ B���s�E��񘈓y ?��&B�u�I<,M���9X �`r�G˧&!7���J�Gɵ�l�cA=����78:9W-�[���1H܆����q-ʖü�O��uv�� ���=�{�E���
��q��;�6!t��ߨ�6�Fe�aqA�&#�*;������I�I�kd��W\ľK��<T��s	$b����u������B#UB ����:
`�`lL����yi��4G��Z����L��1
��e΅��1J�l�+�ᜢ��S�e�U��OXL�K����m��t�uM���u8,�Mr??d�M��s0�Z�T�������Ko�?"�S���������!)�����w�6�7���D�n|V,Y�������w?Pߪ���4F��y�Td��g�Nd���A�˓��6�x^�PӸP_S�DX�]�8v�c�!�����iV�e��2`�y~Δ��9�i��Q�V¡�]1Yiv�Zh���Վe [IB�J�~������i�%K�ZfBz�U�G�^|�5��ݿm�B@��G��4aw�҃�kN�#��M��i@�z��f2t��hrL�������_H�3"��˿��9��;wc@[f��#���p�t�+"�0b����V����{�H�Y����
�;�3ʜ�ϧb��^\�9�b���\��:.�L��Q�@U@PT?y�ī?�ˉ�G{�+�P^f�t\D��m/,��v]�<�9��CЫ�i���8���a��%+��OQжf-$?��qIfmz_�8���N%�؏� �x���P�>���|o �KQ�#ȣ]�B��^��/-�@���T� �.�t�M�#��5�1lBb�u۸�V� bS����e��O�����WN��B��r�G0��������%����;#�,�ǡ�
g^G>������d��b�=���L� �L�?�;Q m@}�����:`G���-[x"�Me��K&�r���0��]�����T������"��=�|�X��-�J��W�Lv���n/��at�>��M���c��X��4����U=��p�E�O����oOG��cL �Z��Н��D=Q�A!����t��r7�{@(���pJ����CwJcm��`��"[��`}�W�>\�%^�dY�q�RTB-W��&���6z��:�Lxl��6"����u���
�'��q��(�w?�Z��U�X�� LR)7�6�4-F!���p�	�W�|̞�P��������?�;@LЌ�g��٭�&�X�ndOH!�"_hGh�����E����^BT{(�5B�8Az�����#���%�ঝ�Rx��Z��8NTN�!ۚ�%3���\�m��`���	>�
�>a��Q���������E��CT���hEhJ2�r �;�,����4�0�x�����Y�}yI������	4�+���;�DGmI���O�H��2�k��O�0��@�a��v+bFP�(>ə���,.��;�u.sd�j��t�$vJ�1&�v���A�-�̊S�С��:H休��jcT[�S5]�D��aL)���_��\%s>:pG�p����=���X�Q�˻?I���	��>�ats �	��*�}m�����ʰl埌�19d��^j��;������tle��WN�ԟ�C�bE,��k�,����5N�R�(���(	�C��-H؟���ڱc�Q�`�z�z ��=Y�z6��>��~�g, ��fzO�/+P����lA�=��P�*}�p�r���>�.�7��'���E�X�C��~]�#1�=X�>,�R/��������Eb<��/�ё�%ֱLT�y�$	�
�ѥmt�h�*�@X�R*�z����};���t1×�xBF�'K1%?>����Ē�:�BߝqŮ���(�����+>;�6�GE��r�D1�Y��t#�����r�k]�u��x�����JՇ}�#3�k��Ԓ.�|�%Uī�����ȥ���~?�a����d�ɍ�,'"X��B�dǠ�Y�_x�W�+w�h���k��-�V�*�j�%��NÃ��z{��ޡ�� P�"�M=� �j���D���o�ODn�(=���PCS;��>���Kw���:59�@�����%��k��ӸY9a �V�R�~���w�y,�8w��̃'\�g�n�fv�kD𰳿ܽ��7�T�5�G��O�����.1�S�m���X9ϧX�Q|�tTq!Z^̳{zQ�Z$`�Ԍ�%��]�?
���S1��k�����2V2RW��]@�`��>��'!��m��$���O-�s��g��q/d���oߘ�E���\m�R���c���xGA�1E�6�3%]��VYƝt��B�W۶]E�2�Iܒ���S{~�q8����ސ�1V�Rz�{�#�-��ͭ��|��BR;@�3��8�\p�h�e���C�F�\<�4�U�~���\7^TN��	�.VSp�!� q�&�$����5	���B�L��,�X �e�$�dY�;����sԆ�Bk�������A4"pyK��<���G�%UqX���y�UX�	�| �ՠ!7nX:�B�f��^��1Z�E��5dI%{��@w��I��of��6�2�G��[�N|jۖ��Y����Jx B�j�Дf�]�x�WByX@`���3QKW����&YRH��J6�,��sL�D_WZ3�:gE͊w
�0ӯ�n4��@
#7�32�R�p�ȴ�B��%-&���t��S�c��<^X�d�&8Z����|�9o:\�[����oj�
rK��gZ��J'��M�^c����v �c(�j�t	kO�� ^�.m�����"}�a.f����pTK��:$��L�-g��N�@Z9M��A���;0b�����}�G��]F:y���h�����|Zt���1���jգ���yl2ꀨ�r5S����`��K�(uzO5�r����ڕ�wd[n������ѯ�����0�e*�N�����%��Km��2���+��4\��k��8��Z5�%����dޑ��фI��^�6�Q��^�o6=
�X�m�I�ٻ����H_�B�Ŝ����_/��G'����+	��a�kAH�H�\��7w�:��Ò �}u�1�/l��n�a���øv�N>�;�yZ?�m	z�΁<��J��ׂ&�oJ����؎G��0X�X�z��Rkf>�e�F�*�)?_SY��c]��
�Z.��N�ѹ@į��(�o܉ X�&hHb�Lv�U�j�m��`Ov�;�_�sѐ~|�T���Std���Ñ�u�-�%5���t�P����P�K�G,���N��#�[[�W�Sfl�aZe@3*��İ�JP	��ٟ��x����w�G�3��ç~^��d�&^���v��V[�����U!��q\�6]���7^M=���+V�248m�M֓N� ��=�׭3'���2�#P�7�ܤ�;��H�Z�xơ�x��}��X�olg���K�����E+�n��E[L8� ��&�}��ژ�y�aK6	�PH�������3P��}�ܖ̓	leQɑhx(��uX3įU��?d����e���ԭ`���2��Scn�{�gSҀ
������_�3F7c�U�LM����Hq����"�\��5� �_�Mp6Q6g�"�L�E�������v������^���fp����E&p#p]���ey�=>������ƴ��÷9lv���*�F����(�s��Ğ��$5��)�le�"ӫ1=��RyU�\OJ	8:���ڢ���{?Q�ͬ@���}�z\�CN���z