XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��o�O���("���{ީY�]IR��fB|/�! 10[l����30'#��V�p��M4��B첅C�\���do`��e'K�)���ب|���G���3a�ҵYA����%^i�玻HS�n�b	��t�}y�)2�8	�)!�M:�@x���k�n�p��d�?�T5���Ȕ�鷎h�z�uϕ�����q(��^����o���n�K�' eX<U�	�����=��k�T�Q�s}W+wo_����E��`�?��rp&�Nt��C�~�t�~۾B�O=�(
�=��x��	��J�jQJ�"b �\�\L���[dpf7��0B%��g�!Yɤ����'Zz����te��Zu�k`iБ��(B�
Җ�d}a�V�X%BXP�A���}�����v5 ��1'C���]�De�	e´�bX;G�wJ=����^0�����=�NEyK,[w�Xţo��l�9�r��j^3��f���3^���y���P�VMGKx�'�_
?������Fw��
��+ܤ�%v��ɸK�x��6�C��6��]/,�����qy�ԭ_���+XNS���$F�|����OTIGh �iX��C�SH�V?yHjT�0����]=I��8棁�Ų	XO?��ܚ=���/���
��� f�T�.?�1oL�0� Qe�ܧd�x8����b����0�$)۸t)e&��V:�\E��M���fAv���3����K�:q�Q8�P\a��.B4�q9!�~�����V��XlxVHYEB    5e2b    1530w���u�?�䁜]BXa�A�#�x�}�Q�2CUa�3�v����Ha#~Ǉ>͏����{ W��.�h=f�%��d¥����Z�o�E�jވړ�(4�qB~��[OTC}�\?�,f��`������Q˜=�KF6�t(`�?�ȑUgD7U��AU 1����+y�opau���ٰ�r%�>B&da��>~G'�1A�Ὅ�o��<���샩K�v��~�BPy�O��yy��
�|��`>G�1���|bͲ�^�Bk5
g�
N���D!�	j�x�Yh�O(�;�	 _���������x/����w�9RP+K����Ep���nX^n�7�9d�e��_�� �f�v nx��ؼ�)�Ԝ�C���6��8pE׌"5�g㾢�j����f���U1'G�G	�"��@K�g5��@㙠��;�;��ۯ�}H$�/�L�'�0�á��`������&��k�@����'ߋS�v����%p��DJOj�	;��{\V�ʫ�[a��9�<C�4m5�V��k��X���)���J[� �:]�_��M}��9r��l�*��r�%O�ت��h|Q�U�P���	?P�,٬��0c6����7��s�\ʄuG��x�3!�#�bi�[�_��Ae��~ǏZh�w�V�����S]VR��ɔ�C}\������^D��aj�7L�@���b繦�`����"uu�^G��8d�R�ߋ:~[��b�?��Qsϧ����c���*�%�ST���z�@����ε��T���{֛]�� �:F 	&�2��"L ��l�8w�2����2��N�Λv4��o�o�~�(�����ɯ��_�1i<��_��|�ݢ��X	Z�j��r��.�C��m���(��}�X��<\v��FL|n�RC���W���Qq:�&,�aɕ��~���˪��!R�ZD�V=�/��̾�q\�>e���0k����s��C7���2�H)���̽���+��Q_\��Ma��em�YB�z?I�Z��bNxȲr;U��W쵐�l>c�Tݪ�%[$�A>MU�/KPu\�ԍ����o'�(�}��d���c�d�����XG������H� 巣�yhMz�<^Ϛ�=�H3��W]�-�WU�,a�����d^S �'ه���<#��p�_SQ�e�m��`�{q~kp����m}=g�{���$�t���O�o�!H82$���w��
ۯ8@��>����^~���pG�O�݉}Z�'����I��6D .?L��B,zr�e� l��!+{y5	Ii�X�tT�uw��p�ǰӛ	��a����)0��Ҥc�����̹ �S�R��Ơ]T۳���@M��2�U\F� �.���C�B��d�4'W�5��V#�a��ĸ���%�e���P��Qv��߷yt���n��p�a�^�zPD����;'V��l�H����	�f����Q�R��P���gz�&Y����'rn;�'�\Sݒx�Q���~�5�'��^eUhN�(�3֜�ہ����H��*�y [0s��.�0�xR��O�/\���� s�W�����G�.7*��9Jc����l{��i��n��\���2E�pB~VS=.�%I;���:�+�A�X��Ӹ�+b�Y�{U/��2�qV_��_]:�m�{x�;֐�xD����#�J9���s�m��򿠥����ԃ��h��(kd��ğ2�)B�ժ@Kw>N;�wAԀ�'�g��CI�S�qO���Ly"ⴑ,���wv�/xr-�b��{�"�z��>�`�S��UN���@D.oj0�>�@�΁�����]Q��!G�"�-��D_�=g>�;v��E��:3e/)��R"�k�\����x5[O�w����c��2fyQ����a ���Y\��*n#�'S��Z���vz�6A�A��Ch��祟(rl���Y���v����?3n.���M���R���\B�2@�T�d�[!��������ʢ�ۖ��V53�!��-Cx�����+:�Q5hwx�a�EN�=���[�(<V��fZ;��+<�xl'�o+?������YA�Py4�O��yy�Y;�Z׌�����M�Ű�A����DCWT�=yN��
�ڤ�fhP���8�K8u�YZ�G7�='-�wy�T7����y(���� ����q~���&��<DEtSƮu���Q:�{�o���2416jMn�s��U #y��{nl*r��<��5��d���ٺq���H	�����$5��	T	jV�M�R��j�'�gW��c%#�g����8���;��j�\<ۀ���Sz6�� '  �a��0w�VU�")�ە5�|� �6Z�Z���;T�w�|��!��B�,E\T�/%r��S�d�F�whO[�G���},�7i=�s�ޣtK�F��׾�hs�>҇��e3�26��j��Z���qDZ�@��>'� ��]ï�|�������3��,�WFw��.�u]a��5`�mȆ[kp��B�3\��6\mf����h��m��?8����f�C�tڹ��k'`���;�M�U�b
�6/�lL����})e���S��~b?��li�n�Kl��޾��P��j�)b�tu�:|�rz�V�*���O�E?���Ok޶`��-�f�ǲ=�>�wg��M#��+o��  ��7��T�sr!�R��0���������*|5w�vJ�c�|�:7X��AԴ�WÙ���aڹ�2�<�B�-��:2n��z�(����B���l�M~ci-�q��zu1�{>��&*έ����3�<Z���R�c3���;�םN~�?�\�Qo���(E"�1��#��������őJs�C$`��P�B����J�����h:NcV<���*9ʓ�2��9Xa-k��  q���yG�	�nC9\#��|ɠCiBvB�sÂG���:�6=Jvcnx�A.�G�e�Q�[|^���	���6�;��c�o��3�-����dK`�(� ���:X�g[O��˼Y��Z���鐽����A���'H��19��v}�6K�ӊO-0�[�����N�A�N��Q��.8�w��\��JAP��A��ĆfRy�'&Y�: ׋�[���Y��6�������K��i@g�b'����\螉)�\�ENӸ�.�� ~�I��Y�;pcʄn>�A�uR�=��q��FB	t�TF^u7��n�P˱��]�u��rK�2{�+9y�w���l���N�ʣ4y�F���%��<������d��	�
��[n��M��@d?�ΦX���m���@:ը��������e0"���]��tM���_0�����=��E݀^�7�'+�L�[�_賧�nD`&	������$�h�A�g�����Ϋ�%���	����^�z]MG�����������!kw���Hjz�"
�O�����L�E��C�C6L�0���}�q�>c[G�h6uy����H3�B��������;�G�'���y�ML��Ę��z��dt�d��Z�a�L5=�<O�7Ye�&��o�<�@^]���q6#�'�����-���Kk���	�MJG��WGx��C�u�|
ٹI��.��Eq_�������y�^�)�p$����l)�2�F͓]�c�����$�T���V��7�����և��`z���ն�\9uku1SM���*;�ߖ�t"�&K�!6�?a���׫n��Xz�^�yj��[Z|���
�P�k��¿�+����ݑ��l�'�7fU���2��wdU���;�gL��RÙ�l�z�'`%U@��g)�Sv��>6'���H�:��q����8<ܼ�b�!�X_2�7��#�������k�Eկ>�g=��$���vD���,f_�z�-O�ҭ�ݿ5^
(0w�	b'�qRr�#.@�7� rMu����G@ҍ��əV�s�0�#�V-𧻓v(S;{��xA�j�[� x�G���M���׽����+�� ��|Q�ʏ�% ���$������g�6�UEV��e�fEO�G�zVG��&T��(�d��>%��)Sʟ!����ۣE,�ۗ3�{�cz�<��.���lWٷ3�Y$�И�1�(8���&��D.3�7��m�HD�����t�'� �V�ް�'�5�6~��$4����Y/��"{���}U��T���JF��&�"WY�SH�"&qt	g��A]�����p��c��aי>�oӮ�=�0x��<�(�6*q��=�,����5�xꭵ�ND(U�q��]�.��3�]"�.s!,ur�,�/�6�]�)��V
D[������J՝G�rP?�=�;��-ҭr4��_
2 �o(��rSL0��8����������-_s5�&��8J�'u���͋y�z~&F.���SV�Mا��ϿUDbN�h�s���|c��=a�)qU�b�-�5�|��p	����� ��~�#�Ǚ���O�$����[e����Q&G�NÔ�/y�,,��
���'F D���J����˅��͋����{����j|��Yrk�^4=�4�rp�N7���4�"�96�1��	�i�|�$'إ|��XK����a�<A����Nnd���z\ǤIf��������h�$_���ȵ[q����*�;�}?��p��j�fnvq���Cn9\8p�����۰t���u���ǹ�hb�>�r��좻9�D�,�N�s��x�&���2�` �����`�䫭[(����t$���7��K>0��zb�CA�C�`��Ju)<,����ɎV���Ff����H��aؾ���N�ً.J�sk;�����T�B!�; �h��t�L��6�����+;����\U2����-��#���-�$U�`u�zH��>^M�`3
�,gy���pZ�Ո2@�ۭ�� 4�j2�p�9��
5m�>͌��v��7���c���������_�.����'�\���x�ʹ����|����Z�a�H{m_]✨��>���������w�T�w�)C3y�s.Y ʥ8�����,�l�BX�C�»�T�F���`Լ��Y[�+{ǦQ�-�Y��.�M7����7�m���fv_[�NY��� ��<�_n�ț�]VQ���1�z
^�A�i^Pt�;�@�n{a*%��<dX����ռ�ƀw�i��]DDy+0��A������o��� ��y���|k�γv��C*_H��]�c�?�Qw~}�aB��M|7�9�h�M�m�9>ǟD8�#�Gd C��Nk�h�y�g����A�����TQ�����6�Q]l?P~rɋ�����?Pj&5����&�=er��zE,��6