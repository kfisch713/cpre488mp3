XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��k'����+� e]��B^q�Q9�����(02����:���%"����򲳅��l�5x�;V���������!���"���1W�	0�-�W�x.P���<��sw�IB�N�oFRٿ��T+�w`Ђ��&�O�ޱ'��E��|V�^�5�x�KA�w]��qIb�������"ּ,%ԋW�V?ٶ�F��uq�>���!���DqJl1�
Vo����?�n�7瑪]����ULΟ��Q��Y�8wR��C-�Ϟo���Ҋ� �|�Ģ�UL��v�ݮ��>�5x�0+�K�"o@؝{7:�[��<���#��!)?�4��0`�ߣ��彑�Ot>@`R�8h��z`�P^ v��S_�=��Ę,�>��y�{�S�^�K��?ܛzO*���=H��4�?�t䰣i�3E\A����0������:aC(+�6�f�/�+/4�*��q�s��"��j�����-��_��;Q�m�l�J�Xg	I8��j2��yZ�0�kp��F�[�Yɲ.�C�N^Ȉ����;WRY��g��4�o��y��^�f�';E�bxޞ"��|Ʋ�O������ʋH&K�{?�/�:�Ũ�ppw+���ԖL^L�^�#%�7J݄��!e����(U��I2�A�v�}���/n`j�|l�FL���v�j�w#�p �`[J �3�^��0뇍.��. �aJ� ��|$�sȔD��\޳d &��:3�J`����A�t�c��߆LD��T����@�����XlxVHYEB    241a     ad0�p�g}�`�m7�K��8��k��SKk�p�U#4�x}O�v[jׇ.n|)2�.a�ި�����A-���������ȷ�v~��z��*�L�j��a�-J�j�[���Ƨ+�GH:��sq�y�Q�0N�r���jƤ"�n$(خ�����
�"��NC;��	-��VQ�L�[xǣ�ʒ�>�_A9��ɩ�:�r\�|q�,A�˵5�5��5d߶��T���tpB��*�(�*ӭѭ_���suԄ:{�8_V�h���7�=?I��T2�*s�	K����.-jiuׂˡ+���/{��)d��9���>'��ģju������P�pA��4-O�����Ѕ's���Erj@��̜�S���"�����S���19�Ύ��j���/&\y��Zeמv��G�~��@��ՌV�c�{&��]\����ɣ��J�/ @8nw|�7BZi��I09rbn�'�Qd��Pxp��T�R�63�2L�fG}��BΆ>��]W�eo�}�q"�f%�W�\��j�F�?�B���Q
�)����H1�=H�h���y�VUܛi�������f#5*��!�+l�1�.@�
�4�1�����n��IK7�A�&m�Z`��W�d��<w��لB�k��e��_���"�*Ԋ�	W�.��,���t7�C_�Ä�/����h�!&�Z� ���ߏ0�,��B�i>-��ʔ�V�&y�n�sf�����F��81Ե�y�&ŎO�+ބ-U�u�s��렗�lv�k����T�T��&hzQ��k�ց3�q."��,WL���E�t��y�S���&unr�(�������G��䡣��EU���+� 2�wb�[�Q�27�Uh���� X�g�\��RY���dL t�F}��8Rq��lw�>2��G$*����I1[0v�H����# ��.�(	�MaF�3���?Yfh�$,x{[A��zȟ��C"��U�2R ����# ��<^]��9���.���č�9���S�*�������|�~p'6<FMY��	+�d�JM�a�|4V���W�7/f`����l�<���X�N���v�Mک���I��j��*fT�F5������mvDT��~�k,��:ф0 ��jp�L�ç���0��~t}(}3ӲS�W����F�G�腞����ǜ�2_b㯫smG������G��O����6�r«ƴ�Ol[�r��c�2�ᖥ��pr�N�Ě�Xx~�����È"<�|�A��H�~W���W�=��ܴ�7�m��U��Sĕ�yn���p���@a`g������ri>x�`�!�����E�Ug���i�tO���*u��.3d��,^��:�(��,��׊���gkȳ��	�O��)��U�L��#d3ͦx��<��(�E����M΀�&~ /�\D����GG)�@p�#�?�aU��zF{��ٯX�ˆ�{��H�QS�L��A��㖨j*X㮶JE��V?U�l��oG��5^L/Q�;�K8�TU'�C}tj�دa�&��c���n��P��-shlsҲ�LNhǅ��$j�����a�+)�\��yN�>E�9�Wjv
j�<�μHp>�Y�#�B�e�m�ʓsj��2�.#�o\8(�Q}�\�q�?�)3$�)gWcG�/��E��)Ѷ%�����u5��HЭ�#t�aĺ�-蕛^ ]�g��\XL<9��K�����n��?n�1�GR0Ԟ-�*�!\s����B7(]ݓY��
u��kNfc�����:�_�5���N������avt��%'ypH1�4	���7�Hc�����B,A����В����f��|�=�A�p�k`��+��eg�ǵw��Ȫ�$,��eUBF�������l� �w*-0J�+瑤o�u�y��\��H,h� �G~�B� 5��� 02��)���Z��Z��,rBeWT�%l}���]!+�(�(z�b!��,ɑ���E�Л2`l	�QU��ؒ�)�Ȯ�P���<g'�댺�U�2AZ\(�F���&�5����D|S5#3�r׬���kz~��:��q������{�L��g�3W��m�n�򑇦at��ؘ�5̴Zǫ"B�x��>�3&O��,<D#{e�Z�]P�zq�b�ط�n/l�Bj��d�/���i�������j�
��I���\xE9����,�4�i]T���9Hj�ы[��2�إّWY�ܯqtT1}���^��%�N�M�j`w��i�_<�{]���xXMO���{��j·*��Zd#�eg��%ϔ������R0z=�R�ĩ܃�|Ǿ�J%��q{D���� ���b��`Xys�> �o�F[��&��B���-$t������!ۀ�F;�ญ��A�����y�c�>��33���õ9 �S5^5]yL>�C��Uה��F�r�1i�.�S��h=���J4��-j���s:2e��'r�[�!7���Yb�`����'�K*�j@=�����^9���w�Y9�0d��x��=j�L�\�V���®�D�a��<0zt��JT������D����*����o�O$Ϛ�A�fu��¿Ws𼕘���n�`Yuu�EE�u�.��U�b��rt3��:'����dS�G_kI��!�Q����X��H�3��r�N��o�C� ��n8x�hj1��F�rmFD#D7G�^���Ũ�WfF���w@‌��v,�F]�z���Ž�����6�	��I�