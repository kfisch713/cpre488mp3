XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����g�ˆ��T�gEp���k�'06l0{�����hic�l���FE�焗�\P�کO-�"� ��R�m�L~ 2�J��رF�b�i���`;��x1(�����/z胜wW1�ܧ�=9�udM�]��i	<+.�"��� G\�1�{�� gf����R��BIR@��}\eƢ�=�C�1X��G�G&�t+a̙�۸*���c����$x$d/�n�T�б��>���Z�GZ��B�������F�&��$7��#8z��=:�fD����@�/���P�9�X�z$�q�cF�r�7�!�N�D�#�N��PC|j1��u�:�vs�#�lJ�^p˳�-�-7>�z�fn$"1�Y6��.ps�Y� m�A�~RV3����$SbmFBA����B&�zv��rҷ��݅��M,���x,��n� ?Cyj��t+z`�'�j%�	r}�� �z�C4J� ^X������v��ԩ�͈��z��)�dn��/�CL���'��RZ����9P=X��F*�M�ﾠ���չ���5֔q+�F��Y�A���}XW�r I���=Ɗ�2Ӎ|Ie&�� �TC�x�0#�m�YB�b��*uvL�jXS���<���5<�(�;�.� ��+-�XG��r{R���D�q1F����M`�l�/c�8V�-���')��'p������.���G�`����?X�)И��Mh�)�-�F&��^O�S�t��w����E+��t᷵��5c��/fJ,VEu��XlxVHYEB    1e3a     a20�' Y�"q
�8�,�9�ڹt��5��ʸ���=��Pf�@������6J�s`�zH�j�t���ނª��kKHZL��IN�d�M��w:>7��,dk�c�,���r�d�^�O71=Ŕdw�;.��m�����S�f'X9^�3V�Զ���Q'���Mc�����g���b��	b�ߒ1M����sayP��"�4[�>���x�����D��t��,Y�a/�$�e?�K�o�B�k����g����ѸcF����v?׭����ØI�o;�8B��n�@QȖ��g�?}��z?W'h`��s�����j����6���o�Nh���� ѸLEF�\���h��lX�$2*q$�i�{�~���
�!b��U�2����]��x�����Y�(�^���l�����2�|եP�nަ��F��f��Ę>7ݥ�x����G�pf�R�a��o)b�t�N�X.ʋ��	3��Iz)��z��Ջ%?,��+���{7!Nf�&9<)���D�)�B�c}	���t��J����b�ܕ����ؾ�wKS����{���آ6o�+f��g�x���o@.���v�̘��p�y`��tj&�Px��2Nng���M͒��?`j6��i�����ρ���1�g!�l�3,*W���>"�#��E)f��	rN�| E�� �t�n�'�	"�g�8�Q��oc��t-��u���"����Y�S܁�0ܔ*�x���D�@�_�{�Q�°�x�:��Rk�ӵ�� ds�$P��|?H�#�<���̳B;9׌Z�a�?u�}X2 ��8v"Aݒ�5��S0|����f�WDp�<M諼F
�~�#�KfR��EO��7��~<t��gD"���[l�&x��c�堓g%b%��y2�ƻހ�k�����p憖�:<9Gi��ų6�r����7��_fP��@����6Yt6W�ohߩ�&7]�V�jF 0H�_��wZ�505�H9�E�lݡ&����l �)�K�w�![�uB��P�e�B�P�Srz�wm7B ҵ=g�kj��12���L�I����� [��0��O �s�آo6AL>�}{I#�W�zW?5~|m�k���2Fߝ�l�`���}u��`^�/�S>����нHM�T�}5F�\i
'-2�n믌�����T��J��o�?��8^{�Id$;ψ���M�GHC��.˱��&N؃m�e#����C��k�"+@������{ٽ~��M6�� S��vi��+0�Y���A��az|'dg��ʬOg�i�ۊdu����:�x�Fd	\�	�(�L�>��Wv��g�U�w�?�	����6;�~��jO��}�@�4��ˉ=nJ�J& ��?���B�٭;�t���-��M�~K��ƾ�F�����c�Y�!��	�8tPO��*��)�04s~m*o"�]�4;�>��_C�b���ta�ֱ)Pme\V�Y��S{v��Y��%ۀz�Ӱ���\�5����iu-����Q�������-&����o$+�D���x����p���F��ⲛ%�����T��O]�׫�R_�y�k�)?��xԯ�󴅇]���w�ĝg�g��;�!4����؋[l��d�y����\OXSLo!a��(�[�fU)��	���l����׽T*�йfB5}��Q*n� y~��$���k�a/���8�}��}�0Ƒ,���X����2N�iJ^�]�o�k3�40��	w�Z��øx���|6h=��F �Q�ԶFo�䞪�mr�H�\U)�T�M\vN�+h�!����3�����sa�Ė�e�B�S��C�U�3��'��2CP���T�V�趟&�]� �N}e�.A`�\��Y �[~��3/R�ԃn�*w-(5>8Դ�ު~H�QƸ�a��s̨��5:��&溍����^]����JO���-��C����N�u�u>������1e獱����+��0$DS&9,��+'M6�+����4!�cL���kgU����7"B+��.v�j�9�R� ��9�	�,��@LT�['��,�;�k���4�ě>-	�(�c�w�AR84O"�#w��ǎŕ���p�3;q�=���+&���~g����[��k!;m��)O��42t�5by�GY���"���Y׏�����A�qb��o�d��ÊJ��6Q�" �?��N/蕡����/X��+�`��l�3�U�:U.���r���}k��/�� (�/*H�jg���Ⱥ�#�BM|�G聤�½b��ay��xCv��;�Yې�m'�y֪ǌVF���It
�����?4�l��po*4�(�mmUiX�Lv��G$_=�h�P	��G=G1�8��b��Ь��J���2��B��:��#�a�� �`�W�Rԭ~��Q����!�6���$�	�V��n�	#��-�����Du�I2��>������O
7" �)�Pr��k,�N��*�X�	�Rj~�M���3�kڛK�q+�+d�z�C(Ŗf���������M
�ٸ{�RmGv5�|���$�k�7d�ϖ�2�b~�忒.V�/U��cA Ҕ��¶�5@