XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�� t���CF p��xwKSp!k2�*��d�4ɶs$��dbC�k���Z�����|d\�jbjxv6�h�ؿ�üU�{�~Vb��Ng�Yn��إHU4�B�������>us|F�+�4+1^�,kw/�^}c�M뛀WK�F�X��Ak��Ew/kV������nf���G�Ϛ3�B�����T �̞��|U ��
�gx����I�w��%�O�\��KV��}���ͻ�������������^� v��\��欺�4e�2LU�&T�lzb�����K�y���F��ԋ(7<wܮ�:.���.�2����kV��w��'�a�5���V}�K[������BW��m����L<���_ٴ���X�V��"��%k��d�1�l�E(���slD�X�M�\�&O���C`��/�\�Z�à?2\\��h 1�!����<y{�N�|��b����L���O��S�1Uc���dE���%Ȳf�Y�Yd����P-�#��hU��^j�hC�=��	��Mx�f.��'�h}s?�KG,D}��G�<�$�@�POΧ����8��`��q��0�0���q@�c��jü��#x��c�ͥ��[C��``އҒO�h3����6�Ir7 �&�3oq`؜�#40���D�2Ǚ���U��2��ڪq-"�l�Pn�*@�I��q Q�rp����C����T'�k:�p)��4�����z��NV�~Ԝ��
 �n��ݦ�'�XlxVHYEB    dd8f    2160�?V�pd�TP�D�Bdb��Nn�� ��*M 5�Q�84qb/�Y�}�8���߽B�+���N-�3���u[T���q57wA�ݢ�A��1O@�sP�����tC���������Nb:��?G�/nb/r�bgw�߃� �$�Vw"���Bۭ++N:�F�ȿ���OЧ�� �n���J���<�yt�׸�t��Y�j?�住��f @��vu/9��R�����s��}��k[��հ�����Ca�=A,����r�Vj@�NĻk7��<X�$�����{s�a�<y����'ɿF�lb�7����O���-b�<�#��Ҕ��FO��u >�<��@z�ɬ�<��������0����J0�$k�\�rdE��3��*Jl;��CH?��3-�%�7O��(�<�pm�uU�=#����;�����_F �-*��b(��JH���Av����;����5h@�|��_�dAp�sX(}F=Kb�,r[�@��/�\qL��k�9�Vٍ�����E\ŶB��몖"�ܹ;����&AϷ����p䭉9$M����o������4�>���s�޾9�/���| �S{�-��#(�p-�/G�R�-�i��h����D���?*�W�,N��\
�	��%�©��$�v��5���Vbk�EF4eS�g��gF�/6��
�P�6-�rZlo�)��y l���h�<�Y�&��Jפ�{�������Nb����x�G��o�uH� �g�R�:̹��������C=�#����]kbd�g��u�2���ܦ�������$_}���i�2��$+�2������TA��d�Y�o{�^��ڴ�>��jw��f�Mo��OH/�?�¡�����ő&+P5���撠2�D��B,�$�J'����ҭ6����墘�+�nC����S�v3
����8ӄ�b��KXT�E_f��>��[�Q�	t"ſGU�y���B_|��%\�����F�_#v`~^"h��N��IE��u���h1����D	W�8p��Oh:%���q�g؍���߽.�=~p�G)���K0)\v 2����F�Q	8T����jOiyh��=���"�	�\��s�!�ĭSa��J#�^��I�P+�ZEe�'��-���U�0i��)��� ��*u�Rzf�Nf�okn�B�u�u.��ZO�ËgEl��8��#K9q�s�w �l�ĉ��f��ܨ:�K��/$�hM^?&�~�1Ȗ���8K�ğl�*<rܒ�~]"��2x��Go>��
Ed��8TA�w;#��b6��9�*ȩg-�i ݸyW���F�s~%�琠~3����K_�;6�XJ�R-z-���H�-̔0",��|El�����F�,�c����5X��	�\����g��]!�Z��-�"�*%�q�i:��!�j�r�����\�(^�q��?�Qot���j�2��V����~���`���-����lA��"��P�&dc��^��DJ(�=���kD��|V�]@�����&J�dhJ�?d�{h:y�K����.��`?�!�8{���Y,�2�)��p�ɦĤ��ߞ�=ѭ]��Qe��FH=�@D��׋.|�Y��h�\Dcr�x�j<G�2�d\�� 2'Ѭ)�J}���6�-���h������Iu�Y��b�}D����4�K��� �U�![S���� tE�q}�/���Z
�[D-��ظ�s��L*1rQ��{	��u�r)�7���#���co->F~�8ұ�*�*�o�(���KP�tf�n2�n�Q�|wq�糰�*xh��:,A��<r��{�Շ�Y�e�`n���������e6\�sP�U�c-�o�7n���Y)�1Yj���bSZH���uQ4@q,��)�Kg����w��~��p�C��Ӥ��z���>3ɡ4�*�;|`E�&�Dp1?3�-�#@�F��'8��y������$�� C�`�ԭ��"t ���k�H�oTR|��	����I̚���O�g:�����&'$"�ͬ��H�艺�喒h�%Q���L�ֻ��`C������`��V�	hWc�K�Sː��l�U�>LU�a��C]���f�v����C�ϳ�37T�s2����>����na��m�{OA�U����8�Q�	�7�oN��0����X�Xh��p�Y%(^��\�1���t��QzB2�ýn�$s�)�M�n�N,�󈕼�:�ӆ.v;�_O<ʜ�0��\�~��QK{O�J����b]I$/�I��L�}���l���Y��V�ڻUC�1�
:#�+�	BeC��d�ܑ�O�Z����`�Ԑ�F$�`:0�d����k��L��	���`��������1�Ӣ���'�p�
��ƙ�Wb��C�7�&I�����E�e,�,�	�f��ϰX����ݡ�n��.�Kl�Ld�l��Knq�q�4N��lD��i�~rD���
=��5���,GŸ/O�O�[�����Hg���۰��0c/���QZ�W/Y��? gm��J�BwEy��~�I^�w��ˮ��S�I�~!3���3Ȗ��(��j��Ҥ�w
lX��@���n���l^��_��@�# ��������@Q6���-#'�֑��[�a4� ��`������,&܋�F�O�����|��)�mMq�n�%��:�Q�>�JT"�r�:�	�	�
_�G�x��au%=�Vt�3�׬�seF/ֆ^��<;��tL��d��}��S�'u��Ȭ�$��y8��כ�h4n'J���W�ս�~E\>�o�~�l-e����(4Ψ
��8UC&۲E�ӏ�J��f���c�x��d�XZ��ͽh{&t~Zb��;�
#������Z�B�f��ܟ���ф��L�7r�fx���[�q	�Uӎ�tr�B��޵5:��O^I�E�c����%�́^q
�Ґ.e�tqs#��"T��<��g�u�e��K�R��,P���tC��YX��zא봜sI)��rr!�դ�@���V��W�����7O��;ڳ3-�u�*7�mm���1Ps�Y�A��T���لh�Rޔ\�WI�*.�5��A.D��]!�nV�6�2ݽ�x"�_JF��C[%a��9�8�
X�c�>T��<a��}Y����Q��b�$n��st���B�����TB!i	̴���[�!v����=a۬o|X~�A�*;�W�j��<�T�m�c���gq��X���$��3���P{��[�ir$Y��,���K0�e��g�G5�{����RO�/�,�R8ȿ�$�S�юe������G7�XMh�+7�d�9p�����O�Z|'`Դ5���0/U����̟�YH����"�m�����g&[y�;�%
������5�爭t*�xV7�չUu`�Cd��4߼���.z�'��W2�R�I��vR���??�L�|4� 2�{>���/����_�BeI2��	���	$�����w6�V�sa�`��_�Ve՞�ni>L��1��Kp���Yw�q%׻P�d(ϭuI����cϭK�)�5C|u3r2.A����Y8%^�e��9�u���>^�������e��j�8���D�j̓�v�ɽ�Y;���N�S�m4Ѹ�t�D�倕�}D%Ϥ�G��ߏ*������![�`�[��Ill�ୄrB<��1��B7�@`8��%R �%w����:vl�ZZT^E�WE��[U�Bb\-ۓCĲm�4>u�2 ��
#nu.])8GR���|��1��v��,�
�'��0v�XqܚS���=�l�� 4Hn]�=K��2��hΫe�,����X�5DR���
�W�$a�NK'�ϑ�<;5�v��!הg�5}�a�A�Å&*�͏�<�\����4[A�~�f;UɅDV��6?�mS�`�2,�;�&�*��r{�B�r����P�
k��͒�����5s��hD5ݮ�\eҚ���V�}6nryK|!W��jn������O Wإ����ھňH���d+5� WSar���6���M�U��g����\S|n�"�Cp���b��s��[~დ��LP��?��]�xg.i>�" sx6!˗)�b��V�l�?�����-vKl["K�H�Ai��k�p���Se��ꒂ4���p��roը3	Gm0�M�n�|������������*��e���O\�d~���Ϯ�A?�8,FZ*�gkʶ\4�#��⎧��[F�	�qXݘE)'B<UX6/M�q��z�e�vOE.h� �ʧ{��7�j?w���U�!�K�?����X���S����}pV�~_�{t���x�L(�1d��DTv�j=���@�����v$��s��5�L^�x���f7�֠�>��~��;��.���	�!�����?_��Ͼӿ���ڇ�"�5�c�)r��w��	ҿ��:�v�}�4x�hpa�ˡY���9yT8�fK�B.�|V��f~n�"�=2Lݬ�T��A�0s03�i85�2`1�t���!�߿�-�VK�H��േ&�bϗ�ϞkAfОw�L�\4�4�e��m�
�����o{�uR�0��W���ѷ�fx����-R%��쪠}�Bh���o�>��_��J����\�/G*�������80�j��)?7�tT{C�8�E�\4^�ww��Uʨ�m�ș�4��>M̓\�c�������,��L漹�*�`I��*9\��I�����]v?Nȃ;P�d����O��};��i�����6J:$Mqi<c#����;A�&���u]��\�*�Ц�|9 �5v��'j�ȥ؊}\���MB.ؒ2L2qt_�(>Ҥx7YQ9p��g�y��P�Lx��v`C�k}�{ v��G���Q��fB$�JxNvHe�P��k2���4%,��B�s�>:X�}�8�e���>�dA!��Ok_IF����{`ꖫ7|�RGYQb=HO� ��.N%0?�%�n�_�6;��DA��4����1h�jQ�'�&rxQ����/�T���$IW>B��/HZ�r`>��U�<׼ڀ��B?�����`�T$l?�i"��e܏ ,8�V-E�p+�L�
�^�����չ�cQ��`�:�>���P�D���=��rL�ɾT�l�hb�����eҙ&���rܱ/e��ڋd��E���_����hy�w�*���Pp|�j�F���߰�o癹F��f  Tẛ��FAB;���y����q���|Z�#�z�GQHz
	��t�� WV�V+�:�����/����{jze2�Q�ω]�u��-C�؄08i��ݦ���RI�-�)Ӄ*�n�ǋ�|��$����|�~\��Q��;�h�V��9��9&��'/�<�:���j�:�ƦQ�#�����Zjwe��g�qޯ�����[�N���x��p�}���� T��P�>�DʁY{K�rK��M����+Z�,O~��i��þz˃2��J��ru����(�y^F[f{*=0�X4`Wn����ɠ������Ҽ�Yz��C�)�~�ͭ��߳ƺ�i�>�j�
s�X,R&�#�}�@(ޢ����@7 �b��X5y���j���G���Gi�K��ed���gy��kK�gj����g��co�Jh0�I!N��c~}���A f�q��x��'J|^-�JT�f�~Zp�b
ͭ��F��\�C���fa�iղP,�*�9!���j&J�F�?ո����ϋQ4�˕�Xe��U;��t�� u���	u:nL}��ު��1Eְ���$�B?g��0V�=c��o(˷�.#&������H��H��a�E�����޹y��&i^V+Yj�y�}���ş������5\o=`Jɋ A���!��,�YxS����
�R �U2�C�٫^	��}U�\��B������s5$Io�_�!ef��D�̦��I:��D	$�S�-/!�{2�?�½^9 ���,�<���1W��V�Qԏvs�*��ke�bw�A2�R�0��4��R�3>c�(�]��K���/�!`5`ߝ�H냻�Ni�+q5��@���X����A~�8��Ф�yvS$��+�:�&�l��z��ٺt��َ�i7�>�eN�ߏ�W�����3��/sc�tt��I��LA�>������'�>66��煽*x�+ID����+���R�m
bj�KkÐЧ�Aoug�F���R<Z�3��J�T�����z��ξ�#T��%+&�崻\�hIa��ޢX�xV�<�ey��*i���fi��`$G�xl�ë
�v9xβ.�|Qb��Tx�J1`5R߸���'�p��u~�[j����5�$�U��$嬯 |_Y��"�}[T[5�*c��^���럕�u��x��Y���2҈ء�/��;�#=	|n#�PM�Q�j�#`�ˊ�a�����z�`�y���;� �{R|��l]�x�9��Q3�����Vb��D:Z�o���s���@� ���w����������2��coZ��f)�@�f��������)�!M_�uN��kX��y�]_����n^Ӓs���7�M�	;	�),��ڨQ���6��(�������1�n�J�M�E\;�ډ��	��]���{�`O��L<�Yo!�l�%�[��$Iy�ֽ62�/%1�/�2:���`�d�߲��N�	�������q7�ėr]Ҍ~�Z;0
S��$!��b�c��� ��]'�Q����4;�V�.wZ#�.��$ ����;ܪ���q��ÿ�^J�j@��P^8LEq���_�*�h���>��v!��0��������l��A��a �qE0��� ����!�ා~�5XOjҎm4W��6�Ł��h������8��$/������;\��-��I�$-��F;+h�<�\Bd`�0�:X�D��HA�T'1S+�'�𷤟+�J����>3�nD��b��}�O��������W�3V,M'���PdFv=¡X����%�Yq%>\>��R�#��gG0�������uq��w��tn5`mP�I�ٛ_Jq�y�ic,qT���2����q5��p�Zf�t|��V���L6O=�Aݴ���PbR�غ���@��}����<tS�)gUG��5X��T��u�J%��j��[���g�*ˈ�|�RX�{��	NA���P��-���a�։��z�韚ԍ�
�ﮝ�c�9��^��O���pGX'�1 �yWBm�/a���cHS�!z�Z���������>����)�%��S�
�5,�X��?wo�^�&�׆4��'�zHE�DL|Нjq���l��<���HW���z�������.�$N
f^��L�R�Ă:����z�I��¼�VܓN�r�b)��gFG�۬���a�ƙ��ne%z�l�U4�;��\:��X$S�><��R��Nr�3߂5����'�o�V�;�*$tR�4�V�������!�u��R�\g��6��q�L��K��<���#z��5{x��5�Y�fӭP�j3�82��7'���}���hwԄ'K+k���S�	��]$���9�Go�a�M1�����s��2�ʎ�3#𰲴�m]Ҧ(Eݳ���|q}�Q��S�rd��Z�a�w��qI:�2;��rS���K�^��Ĩ��b�F�����.��Y�4[�=�4/�5N�F��b̵�XT����5�T��P}n�MW^�����pw)S7�����~vb����c�Ae�����M�d�ahX Qh������'Yt�J�������	����Cq̀��"�x�GՒ"��*�%�A;��jgqk8&ά�䱌�+"-{�Ƃ}����1k�V�W�*Ah\&�G�E�lZ�M'�T��?>�M��{�Q�w��q�g?	i��FִU֣��Q�8a��NX��<�9�'�iAT���Q�A�v^6�W�|�Y�v�R�c�f$x5�p�}��!s�^f'�I:s�ͩC��C��-��̤/�Qa�]eov��V����3�4�c�������fFӏ�2+��I!</�M�W˧�|	A��^�\�&��=�䰆��m��wI�HJ:�����>�!?|Z�%�4�ہ��)�	��])��k�����R]�>Nsm	�O�!��k4�+t|�1y���v�"(="�L��,�fw�?ԷcAUGs�|_��SLF6��jTgS�*��4�p�O��&U�����-^�g�K��&��û��@+��ЍP�v�{��q_p}2�([�W"Cȵ���|��~뇣�M�I_�=�`g���lrޣ�TA�XL���̝�&��X�d�3�������|o\�*_�?s����
����48��7�w�N�Z�Ã�9��j~${�Ñ