XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��4��B7,Lr�Q��*si�_�-�`9:|*�U�K��%f��$�1�{�	˔��a&B	i����_�U���5�e8K��&$�-�D���V8Ca��jn��[�� �χ�/D�@��gO䛚'�q�'�~F`�j�4/|�M�Pm�av]#����+I"���Y�b?��Ո�M}�d���Z[!︥����G,��=���J�u�O����I�����@�ޫ��J�s><��.����N�>��8�w|���H��K���Y�=td��Z]O48s^^��X��kM_?fS���,�|�aT�Gn�ĝ�����Gn�H���Ӟ�x�D�A��K�F����� K32{�*obwr�9C�Ft��d��\T5��U6!�ի�UWD�Һ\h� �]�p*Jz��?�kfDdi>Lw�I���J��B�F�A M��> [��ِ����%�{A`<7��i~���7"�5����X��~�a��D.�:��xf��է���H~6� c0d�"d$#q�`��c����|#��աriHAt$_�m�u�$,��b��I�|�����_z}��P�^3��Qxk,�X/�l͸c��/��� i�Ȁ�u&ʳ�#
y"�#r瓋Po̊?�,���Nw�bg���As���0��E�P��G�)o���)M޵'u��;$�E�^���~�R�3��B[�*�
�%��X<�K�}�Ն��Eo�{�w�_���:�~����g:�,���mx��> ��+�������XlxVHYEB    fa00    2040��(����v� �S>�c|������������TN ��c��cZ%��0����0��� `�V'[jU�3��l'nP�jR
_�|=q�A2�g���c��u9@�JS1�+ѧ��>���esL^����`Ԧ������}Z��r���9�p��P���&j\{4ʋEӡ#���=M�.
VH#�g�����k��dS�>����Y[ٿ?1[�2i`�5ƴV��5���T���D��)缵R_�n��)����36�m��q��e%���9�&ަn�H�N0��O1��dYH{�q�qe�6p�Z4 hx�vO43��Gubdi-'��>��&��j_X�6�b��Cގ{9ttF;�4�k{;��Zq�2=�7٤I�}���}'����ݮ8����͐*	�1Ӈa�s@A��Em���h�6 9Q�	K���P��!dيҹ���۳�ո��B
g�i�b懯�%ՙ��#7��O���gpc�[�����v��f�F�=��lqC퇒���3�)$L/N�1��)��)��G�	�$:�eh��o��	���9��S��(�9�]�I�MiMw���zD���y<.m��Y~딮N��U����yh��=���t�e�V�����x��5�ܛ� �9v:��iJ���)���D�4:l�JΒ��b�=Ak�MNq�8�qYy���t��
!]���\���Y�H�}�~���_yC�<�ӳ��bۈlv���.'yn%:�*%_�		�tt
&\�I�����Vk~ Xke&�j�8�P��a{-�z���A\8.��8.�g�1O��R��nj��0!����}��u�<Ϝ���x���`kt�A��K6�U�=x<�{"oGz�ǈ�|:%*������[��g�j�K��6�� {ފ{�c��De�7�H?�A���a��>?���g�{��'���yA��_7�N���U4׵�����f��lp��f~�EJ�pF�8μ뗸th*��G����5]넰��~��D��/��Ip�z��A�R/V��R��
��@8�lʁ�::( P�n�B�.A�1-�ܡ�
��+�yw�6�U���	���m�o�+_R�P	:�H����m���:�"g�Z��v]�v����r���B?(`��������%'f�'ˌ�'���!XDf�����ׇ�c$n���v�`���8�#T��q����c�ݔ���S�'A�p���7Q��� � ������fjS�!V�Ny�{���!�$g��Kd�����=��O�RD�p�W�w�͗7a7kg��N�j�]\(���!�	�p���"���Y~���}m�u�
��V3�;@�i'�{!�LP�ƳJ�u��EF�#�V�ld���� |��u�&WJ�D��O"8�!K�.��Y�.�4��M������?��?{>C����Ve.�O>�\�$��E�^��D	��t=��q|��.
�j�x���&O�5��o�7?���	؅��;����>���c�W߭[���(��c�M�_���7�����=�l�V�b�"$3{���_��:��>�6�y�M:��u�3���O�l}�#~q�
O��#�`�����5�Anf������}o��\�w�x;��Q�d�Q��F����w�f��
z�?�˜���tN�Rs쯧,�
=�.C�H۽nT�z=�dAm�=6&o���
^� "�/��(�j�����-�C7Ȋ���HR������ �J:��U{�ź����Nk.�ئ�S!_�f �%�%�=�G;�n���)h/_�ȯw���-h�n� Md�Z��o���R#	%�N��1ZCb��J�W�~�4cr�������]4���~�V�2�����x�^V���x��������좄� �ʔ��/�Yٌ�#!!�ފ�lƗע���Ptb�!|1�ص������#	�6��+�w�3BM���<���0��\��5��O��!x�1h_z:��M�J���c<�=O�x��k <*
�n�.e�Z;�m5��}�R3��<�e-I�� x�J%A0HK�z�z�"1̆��M_;�~f���Q�,����;��5��i܍�� ȼ�j�4��y_g�ҩ˄���1�;��n��ۄ��Uv�҉ёֱ���pܤR9y�S-&D7����3G�ӿ�#��
�^p6�I�-W�ώ8(�8?�t}�F(o��U���{��z��3� ��4��Z�|û�|�Uմ}8bП&�1��d�?��עo����Qrꥴ�@���2��t�����g�&�[�<�P+eŉ��9s����ё��Po��D祁�=X$�L9�φ����tw!ia�������e����?rP�d>�|&���2B΋�V����pj��)�ƥ��؆`���w�ÜWQ��s�q�"�H���/���<T�kx�D�þ=g����L����P�[9v(C*���n����:)��K�����Zz4Z��Jb���׺�2�M*�Y��C>���Y��2hC��r�_��D��Q���=frl����WR�M&�Vc��aRwS�������D�ƀ���"��IF��d�N�#ϡ�� f��!.����\"F�l���b<��ה�|C��xj3�.5Y ��E�I7��Ńh���r[��l�box���hr��O�7tX�W{�rb>똑f��[]w��x�j4?��^�FN �7N	Js���^��=���1U����C��j���+����75iJ���U�<g�'M9`�!������<��\,k@���U�$�_���6�w,���ȟh���u�ӟ��X��q����d �'�sx;�Tʂ�l��+4� �X(G���n.qh�Τ��r�@��n(v)?�fP5�JS-k�?M��v�ʆq���N7;?h�w�F�7q̮\a��Wti>6L��Ŷ2��L�wv&�ؠ����uRt�	daB~�i�e(��&���(��2A�|�(,�^�52��*�������yY����J�r��8ӕQIe�/X���I��9գ.�H�Y685��/�]�ڽ�D��[b�L#I��C�Z��*�)	-S;}�_��[�R��I{2�T?\
u�
�)4���>�0� a��|���s�"'g�x�`�(IĴ�t��1�@�։@�:��.��g]tQk[P�|T5I��z�/���(0�f9[�I����%%���g4��qe�|l��L4�,h�{QϹ
y�X޲ISiޛm�S&v�}��Z	����s�QP�ѹ��/�c$���[�>9�j@�t}��m���Ήz/w��ktS９$��2��<������f'����) �]RF�C�w�x�A>ɘP�������,�|UBֺ��	[�܊�l����n�;�S��i=~��11�Voꉒ�����RV�aZrpp|&[����`ǔ�B��Н��m�� ��L����\�����ɮej^�2��r��t�j^��[VS|fs��#�{�A��U����sA�cy�F��S�NY�B»�p���X#�.� ��&u�x�RD�э'�#jZ��p�OTkz��e��@������R��Р�4��3��G!���+	��&-׬���'��L�U1ġff݈���WH���p�e�i���Uj�!�!�&|q`���bT= �(��8K�%�ѹ)���,�Z�GD?�R�D�����KT�k�H(!�G)��5"I"rA� <Y�c!�B�p��5��'M�[+���R�ld�T��
�7+�#Pl�oa�uuyG���<�L�W1���c�cu�dܢ{�:^��$��҈f��6q�$�(S���A���6S(���ғ$zK,�q��������/b�l�qp���C�N�F������:�}�w�"������>����1�4�zN� ����O�s��s[�o�ey�_/^[ۼ�!�5�o�}x{^ಛ���W�[�n˝їK��Z��+�B4�w^C�dZ�����4�9�"�W?E��T��(	w��<�������m,)���9Q:ML;Q\.�á�F ��^r���U����T���$�m�� =��f�F�B�h�^�1��	��O���#qo���^�;*n��a��50�}�X�V[Al6��S�L�l:\�U�n�$��^�i*��f~9��i��<���QM��3�gm�i���+����؍g�7��zd,�`�5�V˩۬$��r9��P��P�t��w@�'���u��(���9���\�;3|�)pE��(�V$e`�R^��-[ŧZ6��"ف5��	���- 9S�V-\�R�J5	KW"*��t� *���԰��y��A:i���Uo{@2�	o>�΍���LۑF�)��Ms���c1��,���[*K�9�S:�l3��-[\si�%K��=���i���g�h5l��;h�?�p�N��3vp9���2;z�w�R�Ɏ��3����9����QX�3��Վ�Fn�K�6�p�Sk[zg����G��a���.���a�U���ٚ�V"B�1��р�}!Ђro��*H�ȅa%f$d@8Z@��3&vQ��_%s�@����	3
��}n�)�O�-z���|����nڥ�|�iS�e�Q6�����D�k��K!�f֣ÀOmI݊��M��7�9k��a�z�⬬�c�sJ+T��I�U&�3[=qDu���zW'ܜ�v��mG�ר�K+�X��:̕��}v�`�!���<��͈� BR'\Qb�_I-�����hF��v���D,u��_#�m�%G۝��޵������Y�zM���~��{<�#6o�L-�h��{��F�[�\�#\%)��a~�����)-�N	R|���w���I�����c��)'�G�!h�q0	$1�R�F��5L��B�3�t��>�dƜj�.۵w}ϻ����m�b
~k#�{��L]�۠-��`Mg���}�l�"�����b�6 A��I/�����"9������z�k���ٕ�����i�M��k�C�Ԟݫ����� ���B�	+���u!�q��No�֯ew������j	�{��P�*�]���=�1���࿛��^1X�64e�m�� �9Gm�ݾ����x�񼽨$����T̯��\����q�ܩ����ؒ�*Ğ�zF����1.<ᗑba7�"�$TsK{lM g�G���
�>Lo�R�~����y!R�I�jR!;ι��G*d��1���pP�u^1\��K��r�x#�%�+P:�ČQ��%qi�
�aٔ/Æ�>'�0���w�qI�Jr��q�&��QHD��!�6J�۫�5��_�����T&�В/�F��rID[�}g@d�ڋg�6��w-���.%��Z!^��]���Y2 ���6�t�;���~/Us���H�E:D��lf)1|/�d��/�q�<ٗ�~�m��;Ŋϧ��T�B��z��U��'��*���!���tʤ6�ݨ�չnd<�_�I��65SL���%��Pk��S>��'��I�v��izl\O<��cC!RA�B�R����|Wg�A�
��8r<������_o���?6 ����w�vo+VS�-uj��_^C�`3+~*�
�4:��m�@y�L�#Pz#��w��v���W�����~�����#(8Y��J�a����C�?;����7ǟB58Rv���u�-���#8�7��T��{5�~�Of����_v4χ����(��"������b���ݩ�#ɟ�E21�{�O�`�c��$:�EB�ӄ�y����v���~d�JbJ�T�Z���u�|��0�L�M�@z����5�HQ.�M��2���n�p)h'��;q��d)�s�dU!,p�3���"��T,u�g�ۅU��o,a��c�	c��*-�H�uS�c�G��S'#{=h����iHtW.��T��I�$�
�zy_�
�q�K�)������_^�n�?��-q*�(]���p�#�dT)C~i	�G8ah��?Ƕ�1���&)�T���fP��u�qG ֥Wp�p.�`8y!�K2�=��U�B��\����q' �}�>�E�SWhìÌ�2�wْ��tc�/�ݎ޶���L��H����^�c~G�{p�J�"�W����/���̶�#[)W>���IjN�G`�q�_���>�q	yN�J�5!o.���N�Yn,,��bT\o��vKr��rtdƕ\����V�;s5v
�f�n �sf�!b��:tؓ�7�WZ�7�ɡ;q{����03�ŀ�C�YDBe������:�WK&9=�|#k�t�!"R��SXٽi�+N;|c�7��r��4��_���`�J��`G�C����r}��H�p5��"8*ːM���)��5*��Z���7g~
:[j��d�bl<+9D�S�I'^���a6�R�H$�c;X��r�._���a���K�G�[�����+<�Y���w\Cm�nbv�g e��[Y�|(u�5	�+��Sv<n�N�4��-1�s�_$�+^:3'%��@0�w�������=P����ǻ���2�Cg� ��o���	���G�a@���������'lA��& ����0߾}�V��Oj�H|����~�F�r���?���FxQh�d�`�^)aM�&	�	��H�W."������<Q'�(d��aG>$I���D؈X�k�H�@ף��k��{��V��D9��$�F�q�˱�^#N�W~�#xUT?7�׈���Y>/�����}b�]�|�i���G���������
AV� �E���/��p*�H��Z �"�#�����Hq��F�$�{�>8�M����۱.����l���=s]�"'��<�[M�˵��I��k��|��Z�pp��&6��Z�~'�=r���iÏ")8j���W�H���u�'��`����w2"�f~��`[<����V4}h=��]�\��N�rn0�e��kS���Zk�z���?�TRVu��9��ϵO��}�%�	;4�����.�g��n��|x��9��l���,���A�a��������m��D�&��o�H2
���	������,i��U����m7{aTi�̰�]�N2�r�Z��u���$���ɭ�4L	g�*Ì_��:�3�=,t��A�jGFP��4��6M-��Y܌��R6��He���!ێ_���I�㚖����Nv����D�V�ҋ��ZJ�P�3
�,\��P�ܣce�&���T���s�ˁ�Nw���>�^zD!@I�c� ����Z�s�}�� MP���ݏ����=��Y�mo~sq�Z�ۃ�`�,��H�����kU`�=뎙�Y袧 �����|�}����ڍKj�t�&_)��G����ST��Et��-���H��r�YѾ+PH�l�q�����x��Ά��M��KGj?��.�B���D)ݗQ}=,����󛁥�[���WP�^i���� �Ǧ���ͻ�j�dM/ yO"*1�Xi*���Z�o0[��f�@q���O�u�_~RN�O�����eA�H�F�I/����8a�l�b�A~qvw���e�.�/W�[;V�L��i2𹖣�����Z}-r�P��r��B�p_dS\��0N�ܼ��n��	��3��&����� �@�7�g��oyq�:n����������-�_�L��t����9;s��׹���o3a�v��~�'�Z4+��A8�K�S;M���,�����#4�1�F��1 V����<�<i̦�ڲ��% ��h��K0����E;s�B��i��'1]!��6�"�����`o.����O�(�fO���Z([>ZQCƜs��\��ؼ]���L��;W�8y��l��)W�� F���E�=M͚k�!�u��A�ҳ}b'*�AZ��s��]�n[���=�m	N�!����bL!�Ga�	����F^[e��s^��)���gn�$�L�	�54��2T���)�ɍmFedppZz����1h�$�� ���b|hk0�*/���p5��s�If�@��/k��cn�9>�|D���<��	��y1B��u��O�n�<H#�6�uY�Av<�o����qȶ��XlxVHYEB    4f62     b50k���f� �6D���髤�7L4�D�W�$�L�Ԑ�W��,��D��G2.?й�͇e�8�hrVZȘ.�����'1@�;q �J�P!c>�n�H9l7��ᴥ�4P:6��ן�+18#��`���ߣ'���� 6�ݜ�jG�����5�z��[T�D$�2���|�5�+L5�0�|�V\�FfO�iо��@� R�'�I��a�$���:��nR
 � �.�o�[��b]w��E�s�C�Y�b��Է�6�W׀!;T�U�mWÐd9~��;U����_V?��nF('�3"YJ|�M$�m˙x�iCN�g7��mɍO�ՏQ>�uќ��?~L����3V�2z�d��\6�Y�	uM0�J'�ds)q�>M�5����s�OR����J&�8�h-�Zt�feJ�.�G�r:-�b"E&��?�o%z�r�s�,����"*�m��ds�����T�lSw�	��-m�aBΦ_����J�E��pr������t:lQx��lVK�o����<3��AOG�"�v�+��$2k��i�ڙN
b����qT7��s��k��`DT}�ض�2�	7���(
A
�U��_/&����� ��l&����J�kŬ+*:ہӱ��\U���&�|	X�7�ӑ��H�ag�j�d�5E��`%<������IzR��I	�Q	���#��]i�񼌏.�}|�#�<��}a���p�ܔ�x�k�4w\��F�	"jr��!\1z���=.<��i(�+���,�>*�7T���ʪ��T�-��J�����yn*�F��Gc��~C�c�qgr۬�(�m�ฤ�>�X�{F��d��,�������Q?�2�T)�.�q�y��˘�cry�z��J���K���@�|ɞ�9l�����p]�����Ox\��uh�L`�nB�� ��P�$�M�#���e��<�{QJ		N����C2�<��n�By3�^�$p���6���Rm�����2�9�'!)�[�d���x�����B
1İ��Ȏe���� ��y����P0�U�d.R7�0�2Xj�z�lc��k����O�.�ӌ�1��\���E�m=�5A�����sUv]d�E5�Ei���]�� ����Eb4��\����#����uR�r���b�Zh9��󴆽ݴL���`Vb��o7>3�e-��L���7�~[�p3AI�jw~ネW�%[�u��][�Mf�a�Y>ĳwt#q[�NR�ٞ�;/zdN�,0-�A訦�!�g(��Q��4;\;�?�� �ѭ�2_�r�Bq���h/�5����{5��"��}�:\�H�8
:$�fV�S��=y��3	.���ϴ����{��>|j�p��K�s��L:;G��d�2��!T�c�j������t&�t��u3J��Ƶ��8�~�I�%q^k���UV3�0��m��QHl�G%�'cK�@߳k�=����t�s�J��!v��WR\�O.vL��M��t�K�D�>���xOCKlf���Q�E�}g�Dy]R�w(����0O���^�^4q=58�z1X��q�bTh�d��m� ��6�T̅�
¼ԑX!�֫�Ù�!��=·�)������mn]4�'��8���6�
>�UƵD�{F���٩ �B�7U�'��їt @��"6�rGUz��l�g:V<�1O��Z g�M�0k%x��L)������ش3N3A�XX�B�/�°�N ����^����֓�����i�����#�\RE��Ȣ_���f�z���P����I�Ji�����@�sp��oAW��_�I�S�T�����AH���O��kZ%�&]b^Ѡ��U>}��y]Q&N#�@.t����c�5Ы�W�x�)l�s2֬.�s��!sv����&ol����y�Ö�q�\_����Cw��hr��|�|!CM	�@U<O��2hKoTn&p+dQ��J)����P����߫�tT�¶c�d�{# Mu��I6Ѵ��������R�
�����{�!���14�1�b�óa���Q��wjۙ\�Cvh�6f_��t�c�X.P�ycV�ӻ�jf�)oC�WM/j��c�Z�5kx��4����J��UJzE��`�;r�?:����  ���8�KY�(8۾��/�v��M�����y��V�`�3j�/��K~�;$���R"��
X��g!��o����[43%���\�5�;����^�	��_q��]@5Z?i���}��3����r]cQ
��v�y�Ǆ�J�N����7�5o��{�8`���^ɓ�.󁬖{�r>U�x�C��\���0h1S���d���Ē��%���J��-�����N�_�+�9H�`�3T9���)L\��e�ϊ���P̎��>��MBğ�f�}j��s`d.{��A��2��?��,������I0V1��]phKgJ(}ϑv���w�/������Ds���L�
O��̩�|s{A!>˞�P��k����u�g8kT����j}{;��
m�г�la�<�{Gʏ��ф�>��Nr<��tzi"��e�H";lto��ZLA��HJs@V0���?�rU"��ls�Ts.�-���,��09Vg�����#J0E�&��L�Ļ�����������IL4K&��Kw1����ǧ�)hU~���ϲ��R/,�A0�j~9�	���q{�W���1s�b�u4��^/�2W��a'<��>��s�ϹץݴU=>7���|H����v�cd:S�JJ��v���O��P��J9���}$�!�%�Q�^WJ߁�K5p��6���W�K0	y��,%���E���L�vA4yk�=��"��0�