XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��N�1�������h��On�R`�[��7�UF�o���vWJ)kE���#h�%�;���&��ڭ�y�� g�AMI	�UE"�4F�"_i�H[nr*�U��}D�t���峈|z6 �6^{�7���UC.��r���GҬv�BDx��%�7�*����#:�)y<3
*��ma��ڋk�O/+������t��D�`brz3�,�EOa�/ji.�%���כ�h4��T$(E��M�L�;@��@���������mpdtd��qW���T1%Y0�sP��*a�``"c��{a��gqqO�|��"]V�ץu��{G��}(����؝k�#��r�4���.)ޟ��-w�ܻimp��/#�S7����f)�F��܅��g������^��g�B�D^������!�*�E��o
�+){���j��z]�1�6��x��d�$���Ȏ��8*S�^����W�h JX���2�ȷ|�W+�J{�%VLN�JSgh ���V����qy��-3�bs�F!:��5+��(6���&�;	��W
�0��]>�9��O!4��N��g�#�-�?pN���C�;f�m_:@~+��}��ι�H;���A�Z��R�j����(��/7�,��{x��k���_f)���L��$���ό %�[��;��(;%�r�+�/!Q��<����{GU��q\�� C��V��d�t�A�7*�k�h��3��T�#C �1�7�	����,Sه�ĵ������$�d-��d' ��DWXlxVHYEB    5fea    1830���/��,7�����)�Mg�P�'5ϥ�Z���l��
�2��|	S��`E�G ���*��٦S?�G�c)�hǦ{��+���ε�t��?�"N��C�2��K
�)�[�u0EZ��]��Pfy
Y��W9'���W�`�{��Ɓ�=��z�eJ��D�j���{$wC�S٦�� zL�+���k�ñ1M�.kr�v�n����b�w�2��x}�����]����Ok��3�~ڹ�/�t���Yp�Z�h��i�W�bl�)f��u�,����.�|#3i�+{6�fdo����L�SL8 �f�9ZzIRbx��?l,���V� V��{{���{�8�A��q�Lg��ف�HgZ��5��	��&̙���V&��41B�~��5�meٸ-��j���d��J�t^�ܭ��	�F;Ko���ĴFO�� ُ���'I���@�?����o��2��L��h�;�v�R���l���}�0���@����y'��}��9us|̃�O�3�����r��â��>C۔N�6�(���X}����:{u~m���U�'*:g�p�
j����l��$��!<A*G�(S���k��5�b�5��>)�]� ���m�0X�/7�$�1�P���cƵ�Iܜ�O�{4H�*��Bx����\�������fܲ8�tk�Cb9��N�(ؼ��DE��I�0�Q9���F���1)�i�J*�) �Q�^�iZ��ߚ��_?EU�C�|)[L�d%�1�N�1����yj������M�>�T''-��v�c�~� ���� #,�9ٌ8M.�WG+v�g�f�ڵ�+'к�]f7x:����oLeY�1�q�L�a_N�|��P�[��=��-���{����Π�KC!hU��A7�)�d�X��4�10��̴�$3Y	Yh��ܣ�	�׋�{�x�؀[2��{R���6b�zˏ�޷Z�)QĹ������8Fˊ�x��G/�����:/� �3��c�����p}`nb�+�K��HjE[���3l9?��D̸��+x{���('� �^�������T{cX�4�w��U��ՂSnP���W��*�� �Ԃj�_��b�:�UUbܵ�:q2>�g	v~�a:֤@�F�Ex̉�_�������5U�ou�x<{�n��\���ܟ|�V�����+!v!ۙ��܇�a@vj�	'�̼��k��S�|.>Qwv����j.HGV��yVp<��ͽ�=�6��Q� 3���Y���ly�T�=K��z������<Ir.|TeW�P;�0\�I �*^�U,*��ګG���eli՘��Q�hԌZ2� �f����b;';&!�Y���A��IpgXyg��r݉X�GO۴�@mЛ3ֶ��B�-d�����Z5���gb�J�9�k�X�{i9<�G!`��XR���3""�U��Z�>�z���'�"��$�Q��r����B��Ƭ�L��i�-�y��ҙ��u�}(7��`�(�,�Т)o�?or�K�U��-ol9l�6�Ժ=�����~���2�A�0A5qF��~ٯ�ea�_�q�Q�A"3�2�CP=_���V�-���z�bj8���r&Y���_�!���wm�x9�n�2;:����hd�Ά
rēl����[�YO���މT��Bw�ʛ�f��"�<I��b�VJyֺ ��h^F�>CΔ���q8��̭�G�N9�!�t���"�&�3��s���D��q1p*�ׁ�z�t��ud�7+���w���V� ��;A��u�ZHH8g��1N�4�xd@4�,�3Vٔ�& UNBK��b榺�jP܁�0�������7�hC��>o������г�@����.&DK���{�o�}�x�I{5�Yw ���!�b�\��N`|���p�|_V!��ȡ���Ff���
;0x6�����j��"���@��24���V!Z奛������s��c�qZ�S�� �1s�3�w��9q�m����V�	R���%�E6�m���U[蟣��zv��7D8�[�� �B��C�<�PD��ٯ�}�6�\��.7�~��;��-8���Pq�_�AP��u���+�t��&c�k�{�721�SȎʰ�L�3G �Q/z�f7��� }sI*� �(���1r�
�m�z�'lGf�x�Ff�t�&Ϩ�É�,���,`�7;K2�sW�Q�'�(�#��Y�ݍ�ր
��+��Ƹ�=��|�B�=�)_ÎJ/ َ��N$�mAN���(\ )p�8���Ǽc��1�3Mw�$;2J����P�e�2δz���Y������γ�������˴���W�E��?��M�x���Mڢ�>�Q�}�!
��(ZѺ����
���tWb���8����a�_��E��\:���4���/�p��Q���r��1P�NyC��E>	(F�o^^ҡ�ǚT0����������Z=7aOw�� �`�R�k�_�	�������ܲ�m @il%Pa~3�g��c���=,&����Z\/�Ξ��Pû,���	�L����>^x�&�{i	5�e�<ˁ�1c4��f^�� �aOM��7������XT=5#���7�w��c���\�=�v˻K�1����U�i�?���@ų9�EEM�3+C�/$�)V��@��ۣ��%�Q4.���I��ǺI]�؋�|�W|���Έ�@B[��4�Du2���=�Ʀ�#ĕ��eK2�~K|=X$-kS9�]�o�f9d�g2�]����
I����KkkAZ�$:��)�t*#�
F���
Z��"T�t:�e�/�H�z��l�{%�)��!Od���4����=�]˷7?��C�G�N���}�8�Գ��=p8\3�O�	< ��L�X�����W�k^��Rѭ����^Amw�gF%b�@X7,�W�����3��Y'��*+1^��]Vm��Xb��w���(�m1.Fq�O���v�&]2#G�iߛ#_5d=M��@M|k=ʌ�c��N�en� �`0�I�`sZ>.���r �^V�6�9c��ۜ
��h���a�#W�\�'KX���.dG��ϣ2 �[̭Z�BFс�ꑔ��+����Y%���b�	�eETy;��n��KGzgf#�wmsVY����Qا��j?���oOѩk�d[��;��C�M��� ����f�X�_iT9(�GӾSܨ[r��&��$�Rִ��U �-�q�`�Y�j�ԟ�` ���6� ]�{��5�)-i���Y#��pjS^̡Z�7Y3 �&���o7he��Z���qC4[Y"Nf$�b\�%������P�p�"f2Ef��{N��q���a����G!vZbA��������7K>��;�ʟ
�Z�Cn����
Ǒ��^��E�$~���!��A�V�n.��6|�]�7��T��.Hj,2L�	�>����y$ղbl�wu��[�I�Qk�E	f+������N$SI�A�*�j��!���x�U���R�u�f}v�9.�P������b�h�:�����k�Z�$F,�g���M��ĉ�/�j��4�D a�m+W{~œ�'$lI�p�0�g�;�GW��qi�.�]2B����҈��?oqN{?�D�\�����J����?��k����Sw�����B�Uj< *,� �Rd�J�!�l{�&穢}р�
L.k8c��P˺�f�P�����J*�k�8f��T�n��r��,�`Ft'l��X-�	�ͯg�nT�@�y�{���æ��mNz�?��j4N���Y�||ϻ�o;�d��1Q�8�[��WO
�������-�z0��J�g�(4(��q��/^�V?��g����	�);!y$j����tvFhzu5�v�*�&Г�p�)'we.�W�	��7*�� 9��/�� ����?L�����*��y�/��g�|Ij~��XiZ:(��X@Y�#����u�J���s��R�;��j^�if��gA(<����-@�[�J�7����2h����=̔��0�gL��|�頁�<r�S3��o(EB��}6�ŕ�s�?���&�	iR=h\5Y��*"�������X��[��EL,GB��v�7��-:�9�6 u�O�ڭmO�Uk��ҷ"�a}��+���G�S��{t��� o�`lIؠi���NF�����n_#C��}���
�e��b�;�#��O�؅��� ނS���E[��z$��"��~��#����z��=Y�K=���W��Nn�~�	P�bX�����J2]G������w��V0�����Nm6���:�����M�	�s�ٺm�49F������,v!|�i&��/9�唪)�N�*��[��B"R��V� B:b��*"�r�ɇXP��ˋ8U�]��7�sW��&��#:v9�}������2>W�#�B�0HY�E\�j< jM���}��Q�q�`�NhLK������{B�����Pu|��  �cC�Q�R����mu^���?w�|NF��!��i�>�y�� ��иE�'��`�=��Ʃ9F�R�>/�	�����t���Vu�a�:�9�ֈ��E\�e����	��eL:�O���.ER��Ɍ�Fi�ϵ�<ǲ��,5w�PQ���wqkW����҃ J�Fz#���g�[��6���;�C��f���.��2~ҽpo�#���7en} ��
Ņu7�{y|��%�����<��2mWr��5%��X���B?c� �2k���E�!Ct$�S"Ġ�$@��|^�T�A�I���dI��D�9U�3/y凖~�#���1V�C���QH���)ax%g}��~�[�O�ΥV?�}�%�S� ʷ�����m9R��e������?�b�n�P�K�eԉ���1}=�G�,;\e �&�t<�D�]�~5!����D�ՙN��;�&�w�L�;�z�c8�W���ۧ"&�Ӟ)��>-�8�����Kr�(�{vm�j��M�@l�A[* �M�7",#�iSX.�-EC��%^#t�n"�[O�n���T��Q��k���ח����$�p2���M�]�� ̘S��2�����)P�"����NڞiՀЬv&������{�B|G����dF�����<#��r�JI������B�zR
 ���b��
}���}֑�~;��4��m�u�wt �j*JKl'7����FD	�7�9ȣ�,%P?;:X��}w	W������/�J|]�T�n
=XL�� 
4+�'nT�o*��$_�.+8�!�%M��|��^h�����$�łS�n���Ց�Z9f��Mq�ꃍ������c�����yu+�7�w*�:� ����}�_1ŭ����W�p��S��YDw5��-��-�"��v{8oy�V@ª��[�Å�Y��}�����qca��h�C�Ĩ��k(��N��� ɛV���X�s{��!�=bRofBw
e�n�!8�h ����9�C����mL�4��C�s�)���&T�5�;˦���x������}�;�E����1	r��	ۜt.�p����J�lRͯ��T
c\�	fd~D�|����B�R+^��B�w�:�N�H1f�Q;d��2G&��#���K�a)K1,V�����`ʡ�UKƲ2L3�̓@�������N��<8������%/�q8=�j-0�^U���Z�#��9iN�_�<?�mrQ��W��S�o��t6n3�Nՠ�H�Ҩ!������I�⌮�e��K{�H)^+��r�^�p����_'����pZ��3�,�/�r��Ӆ<��%�#����2Z�%m��3�GO���L_}�Q'�!���v'J�y��S�
)Nc��d#>�G���2ܜF��.c{���N!�A�B+�D4r #�@U�U��=�~����� �wC��1��I�So�Y��9���c=��~�Z�/��C��M�L����E�bf[��fuJ�qyx�?�=>� �S �g�Qb�7n4'EB�����ã�D�����Lv�_��}�~f�q��x�UTa��&�0�h�� _����W��bȷ��os-_A�U�d��17a3�C������	ћʄ�p+�reA�VĺI�;Ԑ��"�r�ڀ�"��ji��_q$�