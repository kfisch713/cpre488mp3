XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����x���Tk���%mOF�أ�C�S� �QJ��:�۹
*S_�=Ӻ����2�8g[MSu?�US�������'#��u��G x͐/���ץ��PL��B��v��?{�%�=fCO�O&�����H�*����|x�'�bE��U�z8n~)����bI�Ku
\���Y�Wl��u
O�O�i\v�.��K��TF4�e��\(��s�ƻ9�ݫ��iv�&����^�J ��%9{�
�;������۠LjosU�O���X:rqo�6>���ɘ�	����-�N����0�� �fl�O��k�]EO@d�ȥ��"�ݱ�b���'I��������4��(���S��l���W_�T�?[�㟬����N�d�%n\�J���A�J�B�咧�9�������с���O�$���x��Ik��S�}��mI�M�����8*�^I�"���g՝���1n�E8 �7�����d��� �yTL�~*jD3����b�2�J+�ʋ���7ȠK�j%�Q�ۜ}d5������i&��t��R藛�}>�z��뾕E݌_e�Kٯ�����p���C\L���'���N�>;n��a�����r������0���)?i���]K�׳������U'd����
m��o[Ot^�n�7���?.T�.BRŢ��l_u%�� c}Pѽ|��7P�6�Z��6xDL:��6�?���M�!@Ho!�!���--�z��ir���+QĚ=�dXlxVHYEB    4052    10f0?v�9)�k@>7�OP�s�50ĀNo�Pk�� �be�nV4�T�=8p�gg��GAZ�*��^���S[A�ՙ ���+��&ߔ�y��R}��m�DG7��4r�K�k�Pn���!y���:rX���ŴX��� Q#�l���&"���O4e��#��ӾɰѮ��{-u�y�M[,�OK��~+�0Xȸ{�w#=�(¡�g��K1Α0�9ѵ���O�H<�bK��l,Bj8��Aa����Y�@����r{�� ���ȸ�
�&��u��� hK�o��� >A_�'��.<�c�Aw�ǜV;�6�7`�F|*ߘ�'�ڝ��r�ꉹ����O8��G\p����.\���k^��F»���A_�O���;eq��w=v�ak�l�)?Mذ��xـu�(�?�6]�;�NN��죻-����I�x5��Ax�!�&}������)Z��`~���VA�B���Ű*����
w�y�Wd~���`K+J^�ɝ�X������	�-W�r����D� wiU4#�-�!�;��[���U;n��m�3�͌��S��{��W�1��m��H?�`=𔖫�N���۴�	�C�G�)���F�5�t�x��C��3}ͱF�F[@}�����l��d������&�1������TW�W�(�c��w�y8Si�� �g\�aQ��E�Y���
���S,X��G�R����P�W�Y��,����r�$��T�\[L�x��Vm���7�w�{����ʥ�j���1�=H�:��I8p�v�y������64���y�����~�G-T_�s�ш�h��2u �=z���br,�\~8ٱٕs��9Z��=��Ig@C�Ν��<���"	4���o~�P�;@��f|�z9��fJ٬6U0����tr&U�;�lŝ�n�.���v��)&~b`�����#R������F%�����E�393Y��?9�u���uү�"~���H���OC����/�O#j֛Ē�M���)�|�ܫU��R�'$]Ђ��kR���v9�����d���O�=*qIRD��̌--����Ru)�MۊeAhN�H�AU�}�"C���Ɉ<��񨍚�{���OSA�K�
X�S�?rr�G0�uN�!m�>A	gb<�ʅ��E��	L\�5A[���R���5b!d_1#i�gPS�����W���U��D��)X�05��p�scyU���8<Y6�'��|�oS����,:�\�.�o���`�&��C�Bs_S2�@����D��'s�5Ar�~�ð�]����/
}-Џ�;_�#q2m��'�uAM�b/jVN��١���e�HO��Lz6`:�y����N�R@��?�Z�\p_�b�ӱ�]���GK��N��oT�j���#u^�\a��0����L2��}�����v<,qā��\����8�pAݞ�`��[c�Z�;�^������k�3&�k�38&���u3�e�J���*٦�tMV`�������9�T$�}��y����i��G?�����d:}��Ze�#`���Y����TB��0�B�4\��	�[�V��a\#t���T'wWj��^7��JX�M�DePM�c9ǥ��&�5����q�a�����e~���G�$g�Rl�����0��%q��U�O��$�����)ؑU�`&ʖ+p"�yv��F/Qʞ�`��-��Ml~�u�W���t�GQM{�aR�gco_�(<��s��i�i��f�$�34�"bמ{*`U�'|�骂�z�r~6q�,"�b&��N�:(#�w:P��;u��0}=H��&+r�,Id��=Wa#�H�V��Z9����<ǃE�������?B!&��z��7����\���S�#�	�T)���'�R6��vm {#|*'w�V��;HI嘆9�v��J�D�&a�S&��F�u��U�/��7l�Wey�S�WK�Mpo���'��iW�.�����U�����Vo�_��0��Y8�-�����-�fc
�(�O*!�T�g���k��鍇;�pa��[(����>���	�������*�{ց���O�
W�.��8R�vk�f��Xg�C�Ί�+�4���"����T��v�*����T�:���|��X�i،vp�Bu�.��$�왦�0�A�~I����ܵgVȧ�j��v&J�i���"b���b�P@}��9�	�ښz�'�Λ�@�WP���y�a@��~L��b�Z��kP�i��]U�b�w1&�e��I�r��\ơ�w����J�쇼��	A�5ف�i+E�@jHW�$��5�� 4���;2c�C&��Da���}.<��y4��7�R)c(!���A�xk�V��a��UYH�ű|6[���l��}�\|��B��?=�MD�B��<c``˘�)yL�;Iw��.Y���j��N$ye��z'��J����]�4=�I���o2aYdeߕ��	7��>`��9�r�qa���e��{��.x��A��,~k޵��<�]��J-Q1�y|گ�U� `$��b՗��{�M�]u�G�yԾ�#��.�'g1J�7��2A�� ��(�˨����N��[�	��c'�X�:���nJq�#\�SiԵ;�^oR憒�O�3ć$�;D�XO��v˳��m���ӼPlRX:��4o/��T�����t�w�ؓe�ɸٽ]+���o�+80����kk~.gQ��/�c�Ԋr�7`��نE��R��?+e�kw/Cב�C̒�ǣs�D`�Zo�a4����y��>d�>���Q�/��<ń� M��&��#~�:n����� ��W!���Pc�����q�(��w�'��	ev���O�����x�����`I�1Ɓ���吔��[�ψ#�v�╷E��.����B����ϟD�bU U�w�	7�_6Q=��W|b��&�>#��A����Ԁ���(,�|:������s`����q�Ͳ�t�>�������W�*�����Ȇ|�>&l] m�y�V��:�|V�4�g����yʯ�cX�u�_Z�gMH ��� Ot^��p����?�j��/�T0B��m1_ρ,�򸌣$h�U���dD::0΀�Q����Si?�@�ѭl���'y}ny,�^�C�L"{/ZX:�Ί��=CіE1��/�9�����9U}
���ל#_��I�f0���w:/�=��Gzx��#�!�5c��`"��m$Q�z�;�Km�̑�1F��K"X��-���t�O�U�˔r���l�6��B�o�Uz�TA=�����(઄P���I�n"kɠ��
�yk��iŎX{��| ߉���\ю׀�K���N�{�ӻ�ʝ�nE��E���7ɔ�赵�Y�u�ȔBEtk���`��	f����R��k_S��rJ��ƙ�	\��!5��2k%� �8Ag񄶊�4S,�8T�Z-��K?�d��]J�LT �K���y����U8�Gٹ��b70ÙR	��[H}]p'��J������/�RL���ehB�X.1$�衄(dO��5�x�{�"��c���y!k�M�\�����H���ˇ㰪4��h��q؋|-Nq�ې�t�sYt�.)Z�v�/ks��/����������t)�#z���;�v��l#k�˅j�f+���2���ǟD�/S֤��Q9�j�)FY_�a��I�ri91�>2�B�1���o��B��h�xL�i�WѲ&gR��Y�TC<g�H��GN���49��&vS|"�OD4퇝��
 �ю� `�;�DM��!�hb}��h�J�L�r�j�Z.]��Ӛ�< ?<�X��i�_�j�$t_�0���j!+��r0��)daEfY cuiE�{ª���dz~��`�������V�=� �Ŕ{\��Q�z�#G�(��)�j�H�����$a��1�zw�ί=�� �L����v�5��VG>���{B��|DY��Ȩ�t������~�+\�9����43Vi��L�J=Z�@����f�'�h�*UF)H�zo �](���[�63;�6�G���kI�]B�b�*����W�g%�����#���=��GG�HOi�1�k�h���J������$9�4"�1�CZd
�W����e�z
�Y��o௾��/o+�h�s�ֲ�E��0��ӊv2�w�!7�����嶥��%��sjS�*;��Kp"bj��v{9�ܺ^`)��:�u� ��Lq*�B�����KV=��~�rS���>�x�>ؑE�