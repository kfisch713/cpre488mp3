XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����I��|�٩�j�Z+JBW�V�~�C�=s�	��m��bǔЕ�rோҡ�:�H�/�W�#Λ�=/.��m�Fg,�h�f�
��qve�*M��㐨�������N��S{���L(*�,�a�Jb$�;�
�N�45	A�-��9��ԑXCW/r0i*d��8bp�C8fĻ��6ҁ�Q'SUEe4�R�'���~!�ޝ�Ŕ�Ay�ɞ�?f�|�V��̼��tcO7��A�]�qYA�A�HC����O\~ڟ�0��=�Sz����	�E��v
�t�/�3���V������Cɬ4P�d2°�UD�F��֓�H���|N({����c�a�j㒳���Xk��#9_��٩ne.�'�[=7�H>N�̜	�����6��b(��V���qC���/���Z] f;ޯY�i� m��)-��%��E�D�|�4��	k�{�"p>ĉ3�5�����6�TT�mSz����C�l�瘐Y>�}1����:�-�ѽ����Q=�}�q�_��q7����;�7Z���Я{Qj��s�\�3��~��,��I�T���*�
k�r�J�/���Z�Q�m%ڧ��q峟�Eo~"��
�x�?��p�gT �nޗ�|@iFׅ%
�=`ٸ^��0ca���Gd��mH�|Z+��:[O�r��7�МsXo�����Ս�/3^aĜ��G����4�bӖ@�ҕ&�Gƍ#~�Z��F>r���O�����ht�püw���XlxVHYEB    1847     900�$!�LS)@��?�N�A#�X������J�7<d4t]�>4�X��.g�*�PL��51ɉ��p�sM�W-4���U/��=��b������/s�U�����M$��w:��么�0*� �[�[�6��͖'?��N
��rC�B9D��
��7������.��h�H^�*�(0�k�Ħ��JNP) [W(@����b����/�Fչ�slؚM*����W�D.�h(URu�1��Ik'���:�E^�wΟ�,����F=5 }���u��d��X��=�b�ϟ�$�/��hs�Z.3E���qּc�z��@*oRQ�ohl0@�J����{��OI�*���B/�ʪ��R(ې�[b���5�"��R�>����}�RRT�F�w	%���,��ny�5�� 5��@兗�L�D��A�R�Л�y7t/l�N�B5���j^���	L�m(Y�f���g��FN��Ļ��?S������@�
�e\��c�_[�����ѓJ��T����(�4��������_g�Q��Rc�� ���'��.�Kq�g����6��s�2�3��+t6������/Moso�"�r<��)������c�w��a��X�.��ʞn��K >�i��m�0����D��9��I/r-C���!W��s��b)h�zr��;����ޒ2��A�b��"b��L�!A���U�R��5Ɛ���L	:Y�1����5���A���jK�>�]�|I�+w$�2�%�C�W�U��/���a{h�%�P�[C-2�c�7�2nx����2w}���iq���xq�)�������o�Z�
�)�$:���l��T�|�'��Ƭ���V��H	d�}A#֭-� � �ќ�ڥ�g�	��E}Pãe�)�E�G�^��.ch��*�W��QĪ���>��9x �&��|ua&�)�_�Lz1����P�Y�FV��~��O ���|����K���,:�s���؎�4��8Q�P��%�)8Sb�)��Y^H��֐6��}�Fh#�P�Q1n� �Bݿa��k�o���o����䷒�^��u>e9ye�j�Ҵ��=i9��ʵ�P:�dsI;8���ӣ/xYd�ě��=��8�$+<�s;����}�7����з8���s^zm$�S$�3��\���t�ݙ?�˵�(Ҕt�}���Xp�*�:������ +��Om�e|��y�]Ł3M����ޱ��14hS9@n�)�m�p�l�����Ԑ���Mѹ=5S4�w��z~��u����G���eN�࠷4����D�����DA�X�2ĤF�m��J5�����V�����lu�䢥��c�"��n�ЇF�v̭�,�±�s:t5��#�����@s
��|��!9����Y�׎��M�iI\qf��*��}0;̿P��v'���N����}Ԋ�ɫ�u@�?du-ۣE)+��%��~���v��7��#���,zΠ��g�^ ����ի|��WV��^pj؄)���w	Z�u��O!�>����	5�(�+6���Jް� ����%�x���H�B�wa>��73�]�6
׬�F���5����G�9-�����9c�v8�6�d$,�Q����\��!Օ��zM�)#��S���=u�S��m��3S��E�Z�I��J�H��@s4w4׭!�]�-v���N�D�Z{Z#@�~la�}g�P�c�ie��4 d'�s*B�7���A?M7;(�v��h$�X�a՗��o�r��]�u�M��w
�Bq�R�� ;3:��Da����6	�R�R��x�yvSm¤��e�0j��/k���jӊ����)�BLX>���ys����^tG@�IGO�i
^B8T�b��Y��J%!ӯ�l�Ԃ�%�{=kO�+���/�XQt�������;�M��3P�jPn%���#�QD}x#���TF-�ԦF�1r���?��F�d? UY����y��b���pH=��Apm�nWOړ����E�&�u%�E0�Q��de�i�ܡ��X��;�l��A�¢;Tpj�
D-g�%>�B���xM�Y�VV�Z
[t��Ѵ��胝K,2�8��K;��$ꀌI�2R��G��ѧv��If́%k�T �fk�ə�"��?��pCV�����U6Y��FKЕ�Rn]��kZU�?���%�<�|B�m+�5�l�@lqe/��W�4g(cPV�t��'��U���O���\����0�3R�A��P� �a;4u�Ҹ,As��_)�&U,o�nz�F�