XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��v��F��r�"��@��T(�E!]P�Y�	Zv8<zRP��+O�]]��o1�h4L}�r�TP������9[����ֱ�N��O�8ED�z\��.i��:k�O�j\�'Ϸ���� >�ʳ��h�%ܑ^��쮭l?)�26��o�NL;�LB��>�8�y�`
��j��]p�q���-6���Ӝ�#�J��Qh-����%�G�}����&'?���6�a�RC����|�iոH$�ָ����/
6�v}�Tz���o���6�����(`$eo��|&�D���� ��5��?8��sU4<�_b;Y^��"��es��6&�b~a�մ�r�p�a�KnO)3��`IB�MG_kE�*ٻ��=�r�0^I�L�&���SA���2�>�x����g^5��m�_�<"��l:�K(	�@�۲��E�d'���1�Ņ�\�~7�<�~� �6�_��a�������t��ny>̭�fˊ��Jo�����۴�-t~N��y�'�� ~Őr����`&��}��O(G\W�>nk_o�����F}3����{�lT�?K����.��9r����Q���@�g�oV��쪂��k���e\�K�V�ɧF�O���4>}�������ݬWq��<*�o�fp�&�2p�t�f�fH|��罘_]�m}W��z��**o��X�T�Ru#�w��z[Ǳb���$�zF�>K2@��2g ���YT9Vru"���E���֊��e�#t��6V���mk�Q
�(��Z��|Wcx1XlxVHYEB    da59    2e304��2�W���PY�P`��e[6|Զ.O^��J�0�������X�?Vx�Z��>�H��t���	���eS�M:&��,�%��
���HHgW�P�c�N�~�Kq�(0A�A�
�#{8�9I
��&��_O)��Гr��6���|��ܮ��N��C�UƮ,�X]�����?��#���M�`Lj&u��.�Awq����߿�-���Ib}�u�vR8�
�M�E��hh�ǇJ$�D`7Hܟ��x��R�
�a�M94"qFkAv �X�ʡ��b�o7w]��	\�$AϮ��~���� �Y&����\sDë}5�� ߔ'�2�[�%��O����#M��y8R�B52|����-�s^_����`��~�<��0���۾-E�?'C�S�ȟy��̈�H�A{�X�wsH�~ߘ��4�AoÓ�`������,�d�d����n����4���[:����tLĄm�Y]"sjN���?x�9�P�fwb�N��.�kt�G���|�k2��D�ߓ�sM�a��$�ĳ���������X��N�됆�'�yA�b��8p�Ԁh�U�F� .��3��}�ܪưL%�@�I��J+�k;7�YO�f�}�ZQ����P��+є���N ���&�m�i�4�[ЉQ��ᒁ�v���8�{K�F؋�����k�_?g�0�mџ>���-:��oѽ=��T]���7�4���j�A���q^X���@�clR�N�4��J�n�Q����U"���HS��o������z-?\(�=�n�yM��Zf�`�ܹ|�����u�/z8�� ��8Y���2"�ZRa��V�B���sD�
dUb!f_�7L�������/��ubd̫t>�Jݧ��n�����A��%d�7���Q7����������s���4C]� ?ZT|K����m� �FpST ~�iŁzŪ�7	���)�Ng�
�R�E�{���ߞpu�ŷ���H�7#F�[�zi�-�X��`ݨu�G=Qi\��'o*�MF�p�]� �Qn���w㠵Ѓ))��K���s�a�肨D�[��Y _J2����l/��T6�N�́{�nk|I��mQ�R5�v��������"%=iM"�Y	i0���A�n�I���{�<.։��2a�P��b'�k!
ţ� �|��A��J>H<�ВU��#�)���֛�`���a��"�w���)�H��մU��'�k���>��.�o���u����0@iI�R�����❙�c��xqx&GA[�#oXU���=<(s�X����C�|2���hg!	�)+ߗ$r���S�I��@�᭡���~��y���oiḆ)`7�f�.n7�5V)_�V;7�T���x8�K�ȗ��Ss���s�q �z�m7�=� pI�!�� \_��ۂ�����lK�D�Y(x.H����D`�R�6�iقs��}�$���&���d	S������� ��t�H;e�ӌ1�v���t����o�r����V��]0'{����g	��E����&0���*ƛ�S'-��w��c_"+�S����);���=�C;Ӎ����9�/GJ%�Mm��P��M�-M�WЮ�,a����>(�ƈ5�����,p�;3�,#��-YzĨ���z��������bƿ��(��P���<����9�\���;j,27���߀�[{��vq��|����	��X��?���\�� �)�c-E�2*l)\G0n��ϻ2�5ɸ#��7�Y�|���oB1� &(o��:_�PD �V)�$��k6�߱���jQE� 9��~Pg'�x8�ڜuf ��H�$-=����M�V��dM��Eh�Ydx(	̻�؁��R�b:�n�c� fP��݀I?�sCj8O��rg�};q�@�/�e���x�zN��B[�Z���Șk��-L�̐d�.̻�W���.Fr*���mgGl�Y���{�Գ�]认τ��Ϧl;��˃^t�]�c!Y
��������P�~����<`�c�i�h$�B� bl�fѰ�sZ��tp[�-�8�N�*M��`@��.6�n��=����
��.�eڹfC���k`�x���/�|.l'7�8�sx4b�xw��̭��Q~Cq���A"��I���#ɮ���ި�k�q�z^x���2cp���*�$�(�QXKg|i�1��{�C,ٸ8��ݿ�CFc���8���p\����nۗQ���F�IK�sJ�t-��)���푏�A4 "��w�Fe{Z����H�:^�=D���7�7Bש��#����[��7בֿlCU5�0|�B�W2gד���!�ף��.��7�Z� 5Uh.f�O�NK�n�T�w�e*6$r�H�&P	s�5\޺5r��"uٱ2y3f"�rO[�.MXb�A�gI�s�tH4�g�k�N�¸��Ó�J���㙒>��c0i��F0{n�=�&S1��
�pk�>[2�sV=>We����e����� �*���aih!��Ǧ��{���J�V�i}ȥ�8l��]zlk&���\F��.2dx�7��ΫmZ >K]��a}1�4>@�7�:ln�(o�Ҥ��v���2�#�mL��sq�-3���
QY��������/�6�9E��,n���hx&�n��(��+�v���A����`��`P�_�A�]��r���{!���6:`!��a3e,�<�'����W��_�hӄW�*�����d�B��x��Q'O$\%p!U�ϰ*}�#��j<�^��O��OCb@2��a:�Y�)KȖ��H�L�X�N6��U������B��c26k4*�ys������U����RA�n�o� �h��
��V.5N��R��v>���]x�(�G�:N�F�� ����'v AŐ!f�k�$!�����m��,1Ʃ����.���b��,S��$��Ք߇�#�F�3Jp�g�1��v}Aw�Z0���j�)�k��/S���h,V��4�ͶL��y���e��f�CU|�x��0�>p:L�D�p��Ks1���r��͏���'lQm�t�Ri�g�HFFr	%� #(��QZ�^�?�BPk��Rf����_��?k�3hWO��������|��	Eh ޱ\$X��H$��Mc�PmT*��L:3�9�S����U�~%$�[o�ۓ�pŞFѪ���G���M��ي���2E#�I ����P���6Gy����l��Y�����S���49eL�����x��ŉ�^}��#�
If��d�V4
Cjn�G�����PF��Q��n�c(�kVek���(5:)%�'��k���G�)l*���<�1�Y���Χ�t!?����Y"RI�_3��� /7�1ٌ��N;�kU���q |#,=��qy'�A7�R�_��������υXV�%�1�Y�w.N^r4^N7��J=�7�AU��ͺÓ�v���ia
K{�㰢��~hb�ا�T��pN����RX^gl��8$A�
,�YS¾�"��(ľ:#�"�g����!\��w���% �[�Wn�#?$'�N����y̅1���pթIY�Sc����r����cx�k�>�8�/�d��i�6�0�u$���)X��f?��L�����#,y(#U�ۙg%2��Xi1ÁtU���;g��r�c��K&.~}��0����m*�;�) a�l�x����i�{�$�=k�`��#����������P�)�J���6�f�8/�M-�B�_*^l'����b�~��NX�
���cY1ZPl��e�9��? �\���KS2뱭ߪ��D�C9y�I�y�hӕ"Qot5	_cf�t�fp��@`��X�e��l�\��
�f��|��S�="@���m[<`�;����	���:�I���l�7Չ��]�0�#��KHp�=(i�cw�4k����]�uN�*�87�6#���84�x|�Ys��mv�@�}>��Q��G��vE�A��~��.(��i��+}#4�,-��{Y��\�/��y|�n���U"�C+5,����	Z:V�H�bq,I��t�>=��K׋�x��!��.�~��D0o��������,����7�3d�A�e�V��~��$�%3�Rh���8E�ŋ���+]��sd�,d�#:�m�<�b<�b˃�K�\Y)�����v��Z0����A&�|�"��7�t�e� g@!Xˇ<�"�S����t�v������{�Z�m���#x�֐�<�OZ�K����u�%�t�6B���t@�	��I�{�{]��non�b��X���(MvBv�,�n1�6�����ɥ��:*7�*����'W����q*ګ`�=:� �xcM۽���:�%7Z|i���Ch_��2}�EEE�]� ���� ��P���X�FՁ�ֆ� u�'F�q��!�}�|�=�>��V�6؝6�ye�?g�!ң���>���z�i��F^.�h?~_\���F�ŉ��5a6Ș`��v���4I� n��h|=n��%��P� ���m蓖�}\k��v_;��
��c)��I�ŕ�Ca�Q��L4�>�y�/�7!�[4���zY�8	]�@�,�DW��ˤ� G F��v��F�IZ����;�(����&I�+��B�S
����$>;?�R�z���!�O<1� ���J1��s��R�+��F��nҴ�t�����'�9\����k�� ����VeTҷ:A#�� _U/p��"�ȯQ�J��T	��yF����N`�L��w�ب4	��z�ؒ�u�-jhp�����0��4��`��*�4MN��h� ��/dy�R�-`��NE���1�NW��2��	�V��nUƅ0&�M`z�d��r�L3�7㙍�K`5�u'��I�y�qAĥ��/}��};�l7m�.Њ��B0�Q�D~nNVm�������� ���@�9��cGE�����V+�o|����[�7��R��,%rI%��_��]��?j�Nz����G�1���.�=�ѲPɵ����Y���w�6I��p`��䵜�1�Rf����v�ZW��b� q����/$�c6K�|�#j�oA�`�M��}��9z}��]�0jS����9-��뗘�z��	Lq��u���6]h�tC��9�G��c�(ˇ��_��{<�w୷:�P������o?˘5�Ź�K���آ"i�ʮ��ߛ��6�c@�wW�mD�ꆹq(7�rx����<S:CwAN��p�Hm*쵧5�UwrIAH�\U��fd=jr)ٚ��|:��$��:�3��S�FI���e%� �����p[M��)=�(!�K�^^�t���é��p1��B�y�7�ڟ���z�c#²�ln
']G���f�!�Q�r�{(�Hm���U.��#�kӏ��y]��@������YA��A�~������	.��}c>0�6Q.������0�T�z����b��2�VK��0ѵ�e�2��p���fm���$Ət���dWy-3��e�	~߱�5&�����q��#��HjbI_�X� o��p���e�-��^�i��rX���:D��`FpU�el�9Q#О�)w��ʩ�f�#�@��os����eZ�C��)�O��<�k�	�SQ�"2j8�T���~Z{�wl��71�����`I���}1}��z������t�r)�^x_9W�jeg��;�{r�c%8�r7X��7�����t��wv�P�E���p9 R�	����!�g�]�� �f;�M
|&]�_E��E@ e��W��y����D@8SvDOe}����C
�p�u>h[��0I�1<TOqKO�5�������AQ�]h0AT�4�֝�t-�~(=S�VO2���1�M�Y.ⶒ��j3�/Y]���o�ˮ��/� ��+тRS)�i�U=S7i(���i�����'�5v]k�A��[���YK�,T!�0����w��$�.�v΢����fSO�E�J��d�䇌�f����o��Rn^p�\}H9[$�nNC-hd׿�'�6����G&Z*sc�ӷ'���6�����HD�����Uh�#i��O yZ�y&9Z�͖_��(�/g3ʩ�,Pqh� '����$[d��XA� }��F�w6u����.�y8�:��5�`���0��hez������XH%����;,�;�4��U���r����(O~�#+�R�甡� ky�iB�b4HO^>��H�7��YgN_՜���5��$�'�V��}2����z�P��J|(":E6+55���P���7/�$XA�w�fs����O�չ������S�p+�H$_j8�{��W#m�b����p�o�,����L�UQ���A�Y���<���!����K	#l���)��Փ�X���Q��~9���ǊԊFSw;F�K�&��~����pگ}�� �8��Ds��Ǿ*�~��>�5M�Q��Җ��y�����b����z�#<�1{�~�>3�mH8V���f�p���9�*��C���#���ƩiV��'�9�L��-$]�Ќ��/yt�h�0��<]1P����x��V֗i�������D�X�B M��!cC�G��kؙ�{%h�\Y@���D��=�MP��sb ~�ݒ�I����OTف�U��E��ږ��#�ET9xI+��F�NPm�ر��!�qf�N�O����-Y�<���e�)�*Ec}��_�B�Ǘ)��7y�h~G��=/��FK���m�#Jw8J-��q���.n�R��Ve��o?���m��Jޘq`�4�o2���dA9����?�����Y �3"�.�(X�[���Gkv�-������O+#��%�N�2�9TxAJ<d��<E1NJ֞���k��ҍm�����|*���+�gJn ����!԰pI7A�?PS2�w�"�L1�YZ%�͜�Y���oÝ�.���^l�|\"���JS~�dFk9&}��x�>�'�F�ژ��7���3�}F���Ԙ=.�q���!Pt;G�Vt�	�xa�צ)��0|f���Ͳ[�G4_fT_gJ��B�}�'�I2�ǂ�fXf[2g@�)��B`�e����}�?���s��Ia�y`�'PO�UUKS�Q�#�2��Qt�H����T��c�A�%{�O$�pI�k苦�^���ӒH����ϴ���������Z8��}pn�ƅnW����q(����Ƣ)�i4=ݴ\�Z����ES�{9�������.�V$B5�,L���/�^�2�M���ZT�ue�����k)�>a���k����y*�a�iP�T�`�j@/A�_qeɕ�)�;[��ث�#_*]V�ڬ����42U��5�p�ٓ��f8IZo�#
<��s4�<dz�a`M�Οy�������	 �>i
B�|�2&)I����W�;O���ԛ��d�#���3F猰���� �4kY�.�(��%?1���A�^�>�k_�w
P�-����(9; Ґ44q%/�h%"0,��ĉbϼN���8�]"Կ�E�>�;ޡ���Yk{���� ��O=��8l�0:<i<�)�(�5�J-gh�N%b,}�Υ�J�Wvxjʉ�YS��(
�ܧ�����(��2g?1�cuxƻzʜ� �5���
����Ȗ雸��0�~fo����y"�N8�[gē�i����aG�c:�����\u�'�I^�����î���Z���̽��ƾ������j+��f�7|~ߊMsz�����ۜ��J�ά�}U�!j�S�y�Mn#�U�e"���I=��!K����7�˲����g��SCj>��!6���=�y[��3��Q��yjx�\w�������XF�6���ffC��t�0�-�S���p��%�FUR����J*�op�i���6���kJ�QI��h�%���e�Q��k�\��+�+x�F�nq0�J�&_�����aό|=2iXɶ����-@c��ue��ep��õa-�Y�l��J\��]�W�þ�1=�-У�k.GP�q���B�h��x1��&��u����RʇR|TzC�)�#zx�,��Tt��sS��Ih���7ƀ��c��r>��O`���0 I���^D�e"������8XQ�\L1��`�O�I)�U�S��Jw����<�������A�\:�-=�� �x����)�6ң�m�^���n�boO�+��H�S���"E��v���F!f���!�$A���J-<���,�>ƤD���uR�ifJ�:f1u�ͧ~�pUs[��/Z:s�n�ݟMȡ<��)����������aT� �fW�HT�o���m�7s�t~` wHB1p@×�̱Bm�s�{9%����T���Qf�X�O����r0�bau�>��d�Z�`�zy�4c�0�P����U�� q�}��K1���O�B?@��� ծEɽ�R���R#�%6��w1���]
��I-�f��u����r��� 3����m*���J����Vq�P�lR�$��=lP�4y�д��}���?;]�ub5�Kj}��|�vE�)2�/I.�}wZ4�.TCs#{��c3T鎞-���p���|�]e�����V=�ꎟ����Dz=Li�}�oC�߼�x����N��z	6�Kб��BT����A'~9(�ci��2ZT�蕧1cNk��Q�|���=�ؕ*��k�
�����t5�g�`t�,��T/�W#g8��ƞ �VE4�m7��j΃���� ���6Vd�+[@�_��� �2�c�r���0%!�#�,�#������\�q"ٛx|W����-�6�ĴD��T=�U48:�#6k,Z���.Vz��##\
����ا����&�KM��˷2���^?ܭ�i���x����7xP7�-ݜ���A8mѪ�s2��R�;t�E&��IhtǦ��q֭$����;�3c��9���w���8�y,���262���!�l���!�ڙ{Wnl�g3��U
}�|����(� ��-_)��P�pD�m�����^�--��\!$1�rtǛ6e���F����t��rS��U��=Ag����)"�#�'	f��o��]� 
.�d��P+���S�_�.��۝�)3��_'���5�s� �.��A�}�����q��naufSf���~�sr�r]GVO��\������LFp���̵��I�>��h@�f���9h��Ż�b+[��/TV*l����<%hϭ�֓#�NBЕ�,�g��O��Kv�oH��Ss$�:��ġ�i�����C,�g9_�+�1#�Ds,#�L�u7<X�뭽���9V)�7���Ig��Xj�G��_ī�{��-���"?3r���F��+:^]I�ON�M��yR��&]U��Z�.&����9��!�m�$*��ʶz��WC� �]�����z��1 �4 ���(/�_��f=�0�;�T]��f�c �R ����\�p��yQb����9�:��t\-LS~%5J{WK@�O�tlv� 䧹�Sc��N�?�Ȓb���K{ �WF�4mi3�_]H�s�P͒&�F9-��S�1������Ã�:H�^'k8,&}�C���h�'�g[=��N����Gn,��H�q�0�TW'��eK[�����)� Pr��T=t/����>@ﵤ3LG�ѳ}���+�Y3���Ucq������s���ju̇&�z��b�m�^�,��Dm��^`2�G���l,���&'f���b
kp��?p�Saho�yN(۟�N��1�GD�n]�MC���^�Q/Dy�U�B3�/t���W��l�ے,��i0�Q����p�&�����-���I-`|�O�E��U4��٭*�����^t��qm[����~���F�1T�o����H�d���읫�y�������t���)���`;��t]��O.!��?�93r�pP�Zǝ�0�mR�VG4&�8��%�NM��w�:��5,�я�f[z�3���L6���U d�1 �7�MU O��A%0�hY��ڔ����
,P2��q�Dk.9ڃBA�2��L-$��� TN�����^t��@E}��$06)&u\с���|��8%t�'��vpTGs�<�����|.��aK6��]�6p����]��552k� ��u����	�ǧ�@�[]e��VF�O֊0�j��@m(��dt��E$3@�Cv�s{�z���׹��u���wEd�b'����#�e{e"�Hd��1o#=R��=���_�&y�������n���X�7u�_��>��;v���JF0	���8�J���j�c~�C�^�T���[�����fhp���U�Ձ�՛�B�Y����Pm_PK�t�)��#iW^�����Y��k�|��o�ʴ���z��WȳZ�܌'� D8:2`�S�
7/�����&R�ۣK�i���Dju�&�U�*��-8�FXIީrle*'D��Q�B��,XG@��z|��6\O����SB��y�kD�����5Qa���Ň���k})Ր���T(X(֜�[��*a��w�*+���h����i0o�/��?1�S(����*5��2<�_��� ��>��)����X�]�HQ�H��R�K���jۏoR��� �W��v�o��_~��7��ѤAg(�Q�*�U+ԉ��4\��z'nSc�B�	�*ݣ��������˗��t������rm:�P,��'p@���S��ٺ�{5lz}�ұYR�ǭҲ�q�c:�HS�g�y�'�F�9/Z��a�\�-> %�;edϨ�R=O��\d���=G��z�pZ|=��Ѐ.�(�k��[ڢ t�D�O�p9�]�-��s!#�g`�Y:�q�8�@F��� �Q��%5X��M?���c�f�۠ܞ?l�@
/3�7���m�^j�y�� �{]�"5�_��{/aZQ�ҕР��D�cF�����O�>�FX�kԄI�W�!#z�D��Y��:��?�
��˱�n�g[���5�9�U��ah��]�NYc�-���D�}K�r �����X�n���J/8��q@q��g�0g�q*1ȶ����8M�/��찤u�N��D��J�._��f�Ր��U�gHX��}c�Ղ{�㓄KZ3���C(F=�acyo�-�iǮ_���'�葈|�����س� �ʺ�?�ksv�#>!6�0:"���t3u����}�7Zqn�m�aȁR�AA��T��F,=<��܇Cv(�T"�GӕR#�#�6'Z_C�C|X������sWD۲�eЈЕT�P<%��A1o>:������*��Zn
)�ϋ�T��6��������H�����Mq<���,���;�oމ��e�4���X�O��1�˦B���;17�9	�A����`��,������qk�6�wf����*o�!�ȉJC�]���<����>z����yY��a7'��熑�~�]��`�ZVs.�fK4�"ư�c�������	}��c�� �(������I�)
m���B/Ԏ4�ٙ��Vl9�s��g�wNY�9��D�@�+5I<��MQK,�0���;-�^�*C��K0ݥ�8=���fF�'�TB���;}|O^�#P� �tVex�jD�����HGΚ]��}u��Z��䏆��/��a���MǾj��