XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���Dh� �[٘��������F�����A�؀�<N�K���g���){������#^�S`�-��S��[Gyh,��h�1�^\^W˘���K�T���I�m���-������i8�����qH�������gsR�����܊Z����o��7�(���W�J\+��W��L�w� Idm7e@F�3�]��\~�OP�z�O�0���n���:Ӑ��R͖{�a�Xj������^5�S=���Z�%`��lt�V�$# ��C@P�q��3��,l�<܌L��樃�p���敡=�-�*.xW#���)�	K�a���P*��V�(6C�6i�R�4�ϔ�w7�A0מ�|2P�JF0�j6"��^+�C����GgN�����{V�K�-� �#�(El������E�$�������hq��UW�T�hC�2KI)�\v5)��a� o�����_�Z$�3]]�x_�)k�-�;��\�;*~o�ë`��w�(d2�P$�ɓ�&7F���y�����eƟD�����ʼT�R��H�"8����+���6�5�q�*+Lw�!�$����d�<B_;n��8 3(�g�m���,���Uh������|!�$����\��CjD�T-r��WHh�P@W��D��CAu(�혿Hi[Gu�����	y}�au��q�V��r�k�w�,�yǯ$���b�i��6������|���'nY/�f�/e�9�X�:�/�E��L�[L��$�HZsxXlxVHYEB    15b2     890e�B
H�'�l�+���ޫg���	"�/$՝��	���ku�(��	P�N �˳8�_�����\8�:茛����߳Z����5��ל���)�&K8�E���ש�䦨�$������#��4(0��"t>�������x�,[��r���(����>�4�������b�u)vf��p�VCa\���UVE����4��c�! ��`�,����s=|�}dlM��H>�kX�sP���zS����U�!?F��?0;0վ?NI�x@f3�4LD�	������g����*6:����3E =@�?�P�1;�֕+<��'���'=�T�ƈq�o��TP3���A\��+D��ǣq��� �gR��4�vuk��Hc3\F��B��M!a��)8��v�3���;T�u�C0�����+~����#.��++��R{Q(��9���ߨ��m)��Wh�?s�+�!�������v,u��H������`��Wx��9s�=6���\Rs���t�X뱐>�����q���y�4ݒ�>���EX�R��X�=��	z¥�d����2BW�9@}@�;�/@���U���ɻ�n�ז�gm����Nc�[1&��oE�6�+�S�C�(��b��[0���]_�X�#��AI�W�EVR�p#�3-�jP'TCT ɮ��٢����@�����"ͻ.������FC�Lp+y���tIS%�pKu`���A¢lv�����2�Y0\����;�(y�F+�G�;\l#�+|Қd��&�T��w�rܹ�]������S���y�G�P�L��z��5;�g�4k��R1K�O�3R 3	6�DS}����UB@�"5�����!�4�������F�DXL��J�����D��/{�R��@�9�t�0ʫ*aG��>��-_.��b�t��cf�?��Р�>�������IJ�[=����o�!�[����R�|d8fJ�:����!`�8�>�7Y]�\!6z�˯�W�{�>�nju��UT�!������D��(�J��0�ծ�!�^���c��2���ʆ8���J�eh���k��1�u��9p�qE�Ӈ����2��l����%쉭��-�6M�"�M%����Үe2�À��p��/�I�<���g�^vD_�Tl_�#�af�����2����oP��ę��ݬ�\�2��Չ���Fi�4<�pg'V��(J�L���ո�$ڈ���z�5�l�]~��r�K��9F��Ř��#R�U����l膛2�\�&�i6ths=�s�6-�5�������#B^��.<�,(<�u��!)�{�����1�t@�6!�SB�&��ef�{�95v��}�W�R��qx�Ω>o�!�硯�3l�U��:$Ƽ�ὕ��y�u�Q�O�VT�D��*��@:���vw����	x�Ӑ9"��͝��+XjIѸ�(��e@ei,9����4�s�H�OHR��9s�����>Υ
��J·	�(_܋Y�p��B�D:���*@&4)tTӵ&��{Lq��x-��
��R�	������n���ea�V�\�?��#٥ $�w���ߠ��J$�6��:�s�| �pw}�����.d^ �,�%{�����m1���6�d2�1FI���aY����$�;����A[۸BN�ZT�6���"Bb(���F
�^��g9�\��a����m�0d/~uCdAX�&:�7����Q�"f��O�R��]8���;Jh�:X��-�~�����U� F��@q��S���Z�$�	�J1���f�2�NW< ؃L�I��pk�p�]�����:���Ap/�)�����C,h�&�ȉ� U���ı�4$hh� |�$��l�e����XC�j1�:�*�)nU�<z�rV ������/o5L~�R��G��i����������gbjX���j�B���Hlu�/^�,���v��Eg�@޾COl�!��+z4
�p>����n<����?���j�D����א~�	`�o_���Cj�"��4=����X� �J����L,�ݳ��٣��)1w\r�D�&�����l�bq��Le�L�Y�/'�׭��6����,K��������Mo��~���?�&��)Q����A \V�#��t�