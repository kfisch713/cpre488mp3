XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���N��H��	H�-�s�V���U�Q�t�.R
�k�@����ն�q����+�Z#N����`�	�������r/nj��3�4+����1� ��p
�n����i*��z���)�2#1[�3���֭�fzJ��?��G����Z����HɫG���y��˙*�4�:��K٣�[�Lġ6d�Wq:"�d��'���O�A�r̥������vGP�Ԫ�pDT�٧��s�$^��.Xo��A��6>��U�ty4�Q��E+b�V%���Ls�b��)#���Ǵ�\\�`�b�����P�`*�.
�[�
�=�7I�!��mU�A~����:�2f�ii ��7�`�h̥w7�<BL�&[��b�uS���1��DK�w����$���)�ߜ
[r�F]|�)���as� W���ʒ�g *D߅��3��	�����n�07��8u��q����w9x�b�w�����v�� �)�`Uo+��w��s��ټ�,����\�a��Q4����y9����L�M*-�]X�1bza�퐦7�:�U���
�K=&3B:bѝ���	�:Q�B_wh	���;*�u��*�V�ۻ������*S+^��$����Ђ��d0��m��c�y��2Á
�P3ChafiT`0�l8��e�(�z1
[$�Ub�W�э���DY�z_�\A��)*�Q��z�i�R��A��=�" W�藓,B�4�#t޲gDx����9"�4]�E�5~Ԡǵg�!XlxVHYEB    70a6     b90�R���鑜�ɰ�����6_�Y�Љ�f��]y>��'yp(�.��m:OC�T.���@��`}�^�5�m���Ab�g�A�`!Ԗ�V<A�tG!@B���-��i5!���r���h�݈�@0<?��>l�!��Z*��̾E4F�\b��.JH6-9�ǟVh�~x��Svk��X�v�a�X�{�i�j���y]!R�O�q��ޞ�u $y惡Tt�"���{���܁� qƊ8$�����~0>�o�(<�P0~E:�Xz�$g/Rj�A���v�	"����Ĉ^������t"���"S�lj#��xRxLU�����>C#j]�����v.����7~E����@��U׬UOZ=�]h�~M�һT�x��u%:�_�c��Rֲ�ye#W��/0Vlzt y7ޭ��:U��?eMS ����})'Hx�H-8���(�ݢvh/Lu�w���[t�&ߕcˡp
�@#���{��²h���]���ڪ0sj�-�q�E~���%Kt�01��y*��O�o{�${�R�[�
��fBXOOھ�Z����(;f<T3v��n��ZGR����l�����J"w�i�`�5�d���� v�q&'%G��v'��G+��[͓z��(�����*�1��3
U����:m�<�`Q-��M�z�ò��\Mp���O�ׇ���7�3p2��
+=��o�=�k��������S��QJD�Bҍ�1�>7J|ytDv�3L�k���.W��!M�+2�U����ŏJrƌF������oR%��Y�� N�v>lv�1n�c��žji��K����&$�9����˄ѫw�I��r�vS~l�V�N
sVp��<�0���
2�Bd�R�f*�ai���]n`_3w��H)�������9�yz~�>Ϳ >��JA�B��+�������-~�|u��&���l5&�g^��"�.9?h���2g�+b:�tp�U��e�T��^To�Q4ik!�� >��钚�oj�ӟ�^��qSU�ݢ�U���hi"^%h��|Ö��8�`7܌"�E�l`m%5��{R����y���G�Pƙڶ���Q�c}��,~E���4�D�j|�����x��y�;�c��ߌl��f������Z���<��ч��!ç�/ɰ��ow�ui�����p����ެi9��:��X?exK���n�v��r�0�z����5h6��?5�W�T4@FO��3��^+s�.�F]�Z������ҟΫ�T���B�.Va�C�#��=to����/%y5�p/N�G�FZ�@��4"U�埱Oԡ�	[Fa,F!$UǇ�<��
�z30D@��1�/�T������O���M9>��gg�(�<+�7u�;���9Z�e�$U�Z���9���an��%TSDJ�קk>��vqsY-%������5�:�����B�I�΍a��sx�<�C'd2W`�=�<T6�G���JlB���ۋ.�i�rUI�).�dz�T�h�0AxH"�3�]w��=,�KW���*��Q`��/,�ڦQ�q�� %M,<M-~=A�A�*�Ӯql𨷔�=��ې�4�.��5�>6�P�Y��\�����7嫿NL�j-�WO�Ut�)}�vܣ1�eϦ��8!�*�ЗHR=���fq5���(�hBq�`|2S��_oVac�����gI@ض�����$���b���A��b��T�q�e��WAʆ������h������b: ���d����ez����ӌ����Ɂ!2D�m�&��˄$�THw�
;��d;ͱo<��S+��� Z��G|':�_�������&0��j���e�&=��8\��9�r��K�wi	���?���㳉�oP��7�|/��L,�O4���|>~���XA~��������i&nBBk8,�?�|0L��dU�s�#��\�-��h�+*��ö��Y� ����2��r\QO��Ҁ�غ%~w�a��`�<Ӧ#������#����r#��8��3��S&&�^�,����p\��Ztȡ��ٷ�	/Z7H��� �iKt#�S�g]�A|���^L�Jp�}�ka�h[���87Vz��(�dj5"��k(�G�E����<\��T_�!�0~�i�M��ap?�im� �_��7���|��x�a+��s5U;L����W����*M��$U~<�@������g�V�����_�\|3�������k�������H��jf�VE+澉��4�C��ή�(��n�apqT��_L����+��'==�[t����e�p�Z3)��5�]1�p D��
�:�lp�v9�C���jt��D�m������-�y0�	�^���џu�Ů�͗��'��F�@FLF�ZW=y�d��x���`�c�x��;S�{U������j*d[!dd&CiN�c/%�|)��y��^)F,���%��*����'�Cft�P���ҩ���C��^)�����K�I,Nĵ6�̩D^�;9K���nz�� ��cz��_rS ����('w��4�9��Z!*:��ԃ~,�>̜�N���`��4X�[�՞��v�w+/O�U�?�����T��W	$���G�7��MV_��X�΅�#"�|-[)�H�u��˨k Ӻ��/��5�OJE���~�����Q�]N%����`�����+W����]������qm���yڲJT-й[J�&6���|Жju/V��J�UV�,9���=�@��i����e���n�fpD�R��+"�xq�&���X�t����|�u`%�!��4=�Cj��3Z�[��=�*��2|�Mr�\M:���g�GR��[���^0c����;��K�KT����4=+2�\Mg�x��z�9W�-�~�!� �Z�ڴz�+�F��j�h|k�}����2�w�E�,*��F��1�<��?�Y��f �����(