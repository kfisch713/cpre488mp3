XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Q�	�|��)��:O��"v�����[�c��¢��-��"�9�
o�� �s�����Q�fR;�{NqQ��N7�� SZ0�����]�~\��F�������I���y-���؄#��p����D�Z:~~'	�5�o�X� \y~te���'�e���t7M��v9�}��}�����nb`���*5�6ߔT̃�l`3c��h�0����ƲX��D�������L~b��D�v>l�Қhݫ��
̂��e�����P;VX٧n̨��œ�{��/�Wy��EƤ�eH� Ɛ�`���M�^'���؜�`T�X��F��C-�K��f�;xZ�W���9��f���n�����?y�/��N�¯�g���*k�{�80��7�a��ȸBZ��?z)ߺ�J�!FX[��K��{�~������eA�]E���C��b�Q�֓�T���?����C����rV�e��Z�&x$J��̖�RU�N�2or\=2*?퇋(��d���8�V�����P�p��0]�%���\����W��h=���8��
h*�51n�` j���v�ܴ���ɑ^.��G���0z����).Zp�����Y�����Ňׇ��o�5� ������W�F;�qd��!�%!�ȍO� �ƚwj�kq����Gt�hB~�M�]G��|�Y&��^�%��rc�mY��-q4�'��X��;�������0�ta��pAY�K������P}T�0}�~�.�R���נm8K��Q�So�l���$�l�XlxVHYEB    3fdc    1160φ;M�砙�(�tM�(���,jA�j�������4uC��8FpsF��Y )?�Z`|',e��%�D\&��s�݊�tY��I���%թL��e�6���[X��:���w2���q���M�F�`w0�{�$������������Pw/��u��R�P���3�P�/��NZ���8:ʗ����Pl'<��S������9/��KD��@�B�ˤj����n���BFi��� �ښ����O�[�^rCP`
��T�������2��/��/��
^��Mž�~��HטR��W�!D*�7M������-^��l��8�w}П�n��П%��k��u�?�\�͛~T�U��'��� w{�h���k�_ԔI�	_�T�p
������DN�k:��IWU�giZ�+��4���M���`�.��/]j�A0z�� 3�������i~RDp9�V�ijm9n\2���¿rl�W�ץ������l�5��x�F�5�?},��W�`5�*�ICq磽M����U�$��M�@ڊ�ad�������0
ҧX�^=����PL�/(�X��M��5��� {}�vt�fB[$�Y3R�����ؑ�����,n�;҃��h����O��*�W	�T��b�&���q4@o0�:���✐g��q��x�o 7pٺ0Xn|3p�|_��fldk�|	q���_�,K�l�H�6����?H1�%�U�[�M�si�K����t{4QTX��Պ��N�*��$A_a�7WX~KX�8U��u]�"��"�<� Q2w|��7(8&��Hͨ�/9F'n�ϭ=#�]!�VTu�C���L����[m�7��{���O|��o�v��}o�IW�g	M��\���-?S-@����RN�WߩD�|F3ŋ����mBWP���Cm�ذ �q����T�-����62n��֓���s�c��p>�� �ٱC.�7y9Fc9]���6�A��Ω�p��e5�_��/ifl��H�	��.�C��.�uNvD�7tmͲ�C,,��Za|��,d�� Ǧ�	��'�Ey+[������O�	�ZNg��%��ջ��r^sɕ(���	��d�z��э���!ɕ���ČsC��䔛���m��joe�����<M1z1�d=��Z}��%�#-/�~��m�A��@��tY���My��:P�Y�X�~4F\wwS�@ɪ��t��?�c���7	3����!�[1�����~��,��z�Yf慜���J�M�^9+�n�ݪa� �q�;SqF�!$�s���^���<�9�ȍ����z��9�ӯ�V+�	��H̀A�{��������U[�����q}�55���zP��kV�UA�+�x@�i8�'I ����h�������O.�۳5t	'ks���}M)��	�'��I��`~IMw�C���)���GBc	S�x0E�b�"�j�IN��&Y�����S�j�p���}�v��kD�����mȫ�w ^o���4������Y�\M"��}�z6}#���\�e���� <��<e�{燻MV���k���
=&���8��z��.�Gc�4������1C\��Yၧ����,q�>��/�~~>��)���������������6^���wt�Z�d��~x�+2����-�1�$$��Kԑ��\�oTDg�qD!�
9a�q����k�<��NS��sң����aP���K�^F�	jVXQ�@(�jcQ����j����)��Í֚j]���Y['��������~lʠ����6uW�ˍ��S���o�#��� �w����L�4&z�Ġ+�
r52P��cՑ��ӎ�>n�=k�r3�v���%�K5�N��!�:'�Ŗͼ¤��w��^�[��p���=bt1y�4^�dZN7S{ܩ��de��A	����'�.D~��?,�285H���؞:���'������M/=�����z~ǅPɂ�O��m�h��	c�+͍>r�8�%;��朶a�]���Nk�t/ݮ̿�ea�ҰHEA]-�pY�����Qv�+�kS���h��EiݙĮ��=MKD���ۄ�0,�"asЌ��ٌ�A�7)ǳ<JY�\�^��!�"�\��|f�yq�a9�]�q�9O!z�G�R,�����	وV���uXX��E�ʚ	��L)��F�)�7�6U��3�B ��^�t	eL�|����y�%����L���?M)#`ڴͺ�E��e�x,󟷜�[ˏjE:�S3�[�K���)����3��gG�^�vр��54��3��R�qv��!|����PӸ²*<u{��#j���n"��H]h_M���L7�?�e���$�F�q�j��＀6�24�����_�j�(�B�jB������ܷ�ο��񊲚Tk��S�d��.�ڛ�I=���w����דP��P��a/������:�k xzɓ�^=�������Y7r������ J\�lHy���ϊ������؇��{��$@�1&���Ls!���d�w˙0�;��-���*.��x����2�]�]! ���(3�G�U�{�y�����O���n���2�I�	��H`b�ی�
�$,4�B���V9e~�gy/C�϶7d�?�}�\������i���g�>��<o?n�<�����'��t��N�|�����#�1Kw Xr�43�� �=���ط�V\Y�����<E���/7�%��C��w_*�yY�Њ�zT���K&89y��J��p�ܒ���R�ǛA���a��u���Y�[�Iƭ9j���ū6b!W�5rd*�?�@���2X��Wv���cOݕ��i�AfP�e �����E�\��q��A�YS���1�/ev��ҮS�*ŏ��;��>1U�{I���o'�TK�x�X���bQÙ�Z<b�b|����5lx�=�;?�sj�:ā�
���wb�ew���CiT��`}��=�3m�4_��^,��{���V�\k>������ݺ$�+0��3s&��|�d���ݧ��>�j��H:�����Җ��Z��qI�s���m��^H�uvJ��u�W�/���:���Ԡo�jV��t�4T<M��4���tǐ�W��g����Ҫ��1]�j1l#�	ן�
u
�PS��w���~�PYO���AZp��1�����:Q	6�8�i�R9�_\�#Y
�j��]��2>WS�^���_�mo��>�<F������1V��:x�����"���j���[YR�^1��E첌��t�H� �F��}#dc�+͸tOm'�v� ~²�����b�sx�i#)G�k �ڙ}����Ðh@����lF�D��w�X��� ��|z��}`)�,�.��	N χ��b�`���ͼSs� }����M��?p�a��/�<PK�FIk�\v]j������Z�b��R��'��� �1�!����g��R�Vt�8��mܼ���g�5a�Q�v���(3z�L�+}<���D��O3��UCd���+�;u��y���YD!���x����C;��B�Pq�R��Q�d�G!勽����s�2�4��ͤ���89�	��g(aU�~�Ub��q��\�M����P-b��4��v�.�5S��B_�v��m�����pj/*S�kk�̐P2H��]�ALg'��g������!"�J�4cpLB��ҋE�%�z��/��Y�E��!�f(�k.�x��@��
������a���0#l��,5�3�6h3eN���nu�:�l��1�
K��'=
��/G�5��=�Q���QY�^�~��Ǐw���V�ԽQi�3
Z�q^dg����� �Y�i�녴Э�����`�@��$zT��%�v�皋;7W}0����LN:ɊAI��R����7���^|�ٸ]ʒ�6�^M2��>���e1���$eߊVL l��t�}fqu4��t��P��>fd�hN��g�+���ڦwt ���L0^~�������K���D��b����JKm��,��Ug��M��U���٪y{��pӡC,�$ӆ�@����duP�-ܪ;����gn?v����l^�����_C[�q�2�
kU$ie�v�'�`c���
���K�Blo_����T����ڈ�CO�[6yN�z*�
YL�������#A'�GM~K`4d���|���J-8vI�H�s �.|/��u��ҝ���[�*�1&�����6f<�IN��a�r!��C�,W��i��`�np�o쫼A�˩6��/c��Z+F��`�?���B���q�<��҉� F~�;����#ֿېo�Z�6Ρ���Fq�\.��pw̿ܗӀ�����3x��$V�ټ�A�k���&S*��Ď���X����k$