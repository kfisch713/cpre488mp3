XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��W �ሔ������"���8o�N<�\�%�Pj�X�X���Cw��΅͕\O���+��pBi�:,pm����}YB;�ۻ��ү�iԥZP���@0���7����*�fD���!���0��TiQCz�廅�U����lj�u�jSQ�4���UR[^;�Ƈ$R�Ҕ�M�������,d��"<�+�������_���]D�l:z���'U�3��#\w&rR��붽�2Pp|�`Z�($�v��D<�o��;9�A#��ZSa+Ւ��o�ǂx9
��x?����ŀ�,�En.ȯGv�x�~��z�ڕ�ʡ�}�L�p���׎�K��c
Ui�����^w\J\j"-v�=y�{��B�8/8���2��V&��@:u��e�/p���W��8Q���?8�(�tLT�����S�T���|���}ؒ�JȽ]��kc��a=C��%�a��M�f�3l���c2�v��@$_W��崚Iw#�9��ϭ��|���0�i��������0���D&�>���a�����؜-��?��
>�݈�`r��&a5 ����K��$6L=�i9$A�M�c����h!0��%Ԣ����JrI��GCtJ�Ш�,�-��a*ىc*��?�����O�y����D �1�����Qz�CO\E�����*t�9�"�������r���1¼J�K��E�'�_	�K�bCŐ���kb���l�E�Z⊵g��c��v{���]G_���pL�\=; ����y�XlxVHYEB    15bf     890���1�?�ŧP�d�)�y:��B�VX��{�\�'e�7�m�v�3j��Ju&�#�O���Ǜ�`�"�X*��J}�mQ)���#����(k+g�����}�9�vd�_�'����0�	�yxT(�ۃ�Vt�uWW��.D��3�qhN��1Gč
? %�5ߡ���B���A��\^lk�]w��.�i5s��������c���ց�ں�N��lH~�c�z82�}Ixg��n��"?�Xs�_DBbP��_Kj"�La��~�U��sY�����J'@j�&���!u��!6.\�����O��-���F�t��4��E��-?���([35n���&b"��i�a3�7�%ϻ�������S�k羂d�
�tH��WW��)ޯ��3þ��f�j���0T���)�Q��0���é*��c�O��.n�����H��rj�;���R���<V����-���fG�ܐVIӅ@���ӂ�s4�ZS�!2��g+�&������N��4`�CHZ6a|˃�#8��gcR"�GF����������۾��Z�9�'V�&�^��B�S��xm�j��|�ፇ"q��g�,�"^$����h)���:��^{@����Qg�^wz�L������8���tT`Xf|�C����S��b�Y��XQK�SxM���-��6�m�{�fu���x��o1́{Z/@���"�ý_�1$g~��>VA�{��@62��j,���4��@��Nb+T�ѥ7�E�s��|\�rWyJ�h��	̈́le/o�E~�}��7��+J�<Z�tT�:W����IJEVJ����s��d�oO�h��/X��Z�u�LD�ˠ<^���Y�$��C��#x�N���׵2`#p�������~�ZA)���˲6@Ӝ{#�҉��<J��L�{vɐ��\��	����D|;/]��g&V��[pp!��hQ���35% 2.�"�Rk��@��>��ѣ�Ba�e��M���X�����A���Y kME�I[���-y� �	ٗ��xL�u�B�ZtJ1��í(r׉�St�+�a[����K�g��鞑K!���.��	y��vѡ�RF2)�m������{�W.�/���b��EZ��P=M����ɋK�CSs�?�lݢ�x,ZW��B�X�R����M�1d���VcE�Q����B�0�xˇ-HHy� ��]x��pY�N�XA�)�����۩��í���3/|�#��yd��ho��o}�R����(�~���R����hjGږ�X#�G};"]=�* �CIo~�:΄���Ohd䘱�u���(�����2�d���������՘@�<VT`�(���#�v[j?޼@��zН�h^LN��o`^�i|"*�P{��]r���>����!�C	�N{�2]"@��KR
�h���k~/\���S��\��|yۯ��SQEy\Qs�1��e�D�.��92V�B�bְ�'��̎�y*��l��#���0����l�D�?�p&��O;�k[U��ԂS�?��0Ϩgu2�_`���k�r������!;hJ)n'Xç��ɼ3�85BC�b�5�6�@�$�D��A����v�}\|i�,Wp�e��p��!4�������&����;�DE�5�y��<|A�w}����� ?E���nR��
	�>\Y,��U�W��c����c{��f��j�m�ML�6P�س%KA��F�ԀF�����w�[Fm���W��t=1-�F�v��-�cbcˆF>f�\/:�+V?��Ӛ�b����cp~�0��v�o'{I����_�A�B\U���k���!�_M
��sB.Ӭź�ԊM@���@F�)mZ��(�cEH���Su��KP]�2>^(Fn��H�>v�N��0����NjK܁�kĬ���5�L�m�K[���l��	sB�bf�Y-�߼<�PN�2�����Q#����_
Tjӭ�@��bێ�#�8#ü�i-�Wk�L+���{�����Y���NX(��4`�b]�N��s})N�OS��
YAՖ7�}w'���zb.rH����&��sE�8��S�C�ѥ��򣗴|'��%���gr0K��T�F���0Mtg��*��I!h��
_�ѱTT�*E{�4e��_�Q%�a��a5�r��5