XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���y;3gu#%����o(A&�B�a��Ǆ�SɌ��c�
����
�b��.��Y�hK[���Q�HO��ƻ�"nԹ2�E��b|'�,��A����N���we|�wXqz�TY>���yev�� �+����As	�m�[j4ϒ#�P�����7�v�G�02�������w�.�A�$��6O�(#Z�栯�20�w�����8��^��K��'cX��<����8����\ �l�g#�������+�
�eڸlsMQlE��R&J�ϡ�1�cil{����Ƣ?Fپ�tn_}]�i��.���`ty����J�I�:u��M]��aE����T|�PG�y��� �gC�]ͲI�Q&*�F%�j�����T>Ս�{��Aq��j�Hj��HM�e�Tj��-$�(k��1��GD:2V���V�J1�X	O1Q\��k%�D�������w���]l����7��*�M��1�"���>�3[u?�FHdb��abG��t
����"ڤ*���T�����|�" �t\W#�r�;~��_�oS��\�`���;�{�r��uce�F�*�tϩ�<Pg����j
�C���q���aW8X4�~�lB�Ӟ�,��s[͕r 'M�AJ[E�_�+���f.Շ����8��e����M����q�0��A��ux��3�M^�CL�м�ģ��	�,�����+%H}!�@z$���{M�������R�~�Tkt".��
���߁�RXlxVHYEB    76a7    17c0�K�}��� �ޏ��#oC��配�ۜ�Ӕg&J}׶���l-c"<H'�;�F�{eA]��݄���'��K}^���Z�$r�����v݌��B��=�:O�����$�
�g��D�hC���D�)��u򚩬r����/7۵u�Χ\�KF���.�z+��>���5��	@ ӫ�����M����!��`��Fk������~0�COn�\���/3A1�(��<NChAPR)�Q��vp�G��*�u��/���P'p�A��vtU$mԫ}T��c�(�ð���HU>3%�![`��[����뵏��ё����M'v���c��[��z� L�;f���Z艃>bF-���E�۔�^n�|êi��Rt\ݵwϾI˹�'����5�q?�a�
q�`�6�4$f�\�<ѳ-Ɵ,�ou*��wjz𭓭��=��#������W��rͦ���l�θ�U*��A�q�HJ]�}&��
���-R��*Ɔ7���3g�ɧ����Y����<(��jB��QlýD�ˮH�G�$�9/��{�
��d�kv�܀F�c�St��F��o-��ǈ��Ws�M�>x2�����^�����0�of�b��rѬ�(�A �Y���.�Y{`)����<�)h/t
f���uog���忛^�J���jB��p �|^�#�G����%�IK����l�1�;GsV$���[��d�r�M �
�l�"���G{��g�Ur\C�N�MiIz�r����G������<9]7A,�=�GF;K�ne��&�B��0ǔ �n�t�,(ulՅ�5�$o� ��C���V�جH�|�&蓴j��0F�T�Tz����ļM��2��Gѭd�8`��mr�^m�9��G��O����F�r 5	�m���k(s\�z�{{�r�uY�]KG:o���f/a��V�Zs�	�G^|�Aj���a��j�y�6	<ɚ��.�G�oV�f��&9���J��9�h-�;��PwcO�= �xhA�|��h��l�I���
��.�͝^�^u�Q߫�WLN@#'�2I�ƫ$��6GasV���1:�lP�i��C�����x����Ai'#s9n#*�X��5��;m����(=�I,�Y_�<��FZ��s���%F�>*��	�@�a��w�݀���)'�1�b��1��̸�/�t�9�!�Q�!uS"w�Z0L��5�v|�)%Zf�k(�A��lQ��^Iv��#p�w(�JI��A�?�iaѝ��ct�`-����Ɯ�mh��{p��[k��e�v+��>౼b��	��:`�Y�]���\|5��b�����Y+�3�v�.�R5l���qh�_:��13.c�6��f]�|myq=�Q֧�pq�R�������|����è�����[|���Rw]���4��mD����8ID����BvuL����dJV�w.��*aa��@���)y������wi8M�L�%�����W�� �{嵆�X�'}@`=�[���Ͻ{���Y�F�k���OJ����"(:@B�P4���d^Z_a'��ޭȫe���|�1�<6/��
#h�hx����V�n�.���Ľ�x���5[L{�{Ӽ�X{C!�!�J��}-�6+�~hI]:-��j��[���X_Y��Gwf��$����T��=R�<����r�A�����S͸�|�!�t����á�ԸI9���T�[�f�?o~�~r2BϷ����Y����1�{��X<f�������%�$ƨ�9]Ij���a�|�@��y��n��)e[d���%f!��h]��Q�j�,�S��G�����;����&��$���ESV�;�Ki�[��&Wq�Ca�M֬j�2�T����E�2���J�[nL��2
���k@d��_�c j�5N)K�7*�<IV�>P|��B��"�O�N?%�Wi\��g��z'����m���u/��	|���퐬�O �M�D����s���B�W�}�"�����0f��  y���oD!I]B�Z�Y��6���b����|�@^4�u$���͖Ї�Bю�KM��m&_�l}�a�?;�ohB�xT}L��)T�<��j�KE��r�� �j~u�:*PL�\~��զ�4�F/��E��{9*Nl���#W.9&Ԧ"�c�ݠ9�����J>|�G��nOC1�#���}�f��Dno���P��m�
��Lô�h�je�J@ʛd���2�����I_xש(v7�RŽF�NO�F���'}��j�h��+]��P�5�0Nr*I	�%2ڮg}�����h��$��%��Q	���j]�����yRZ����h�rM�I�����9 |�G�ԝrv�}����w)fT�m�kf�����o��vZ.:Z����.~yyϗ����"�Yt�D����?�D6�nWp��UCn���o����\d����/J���P�*`�^�Y�m�颎��m����K���ZΫo���=�Hp��:�M��I��2Cܩ�_ aD���o��
�i����>^�mf�;�1�zF1�������D)i��3�J�ܔ�]��Q���6��4����43�Wl�	��A#������$�Ug�$�|�p����>�7�ڎ�p�<P��2���-ު�cw~G>o�iDr����/�6��Q��b���SL�C#���PN�%�kSB������L���ly@�z>�4��d;�� �>�0�V]JtS�;�+���3F	z�h������6b�ZӼ?�/(�4��j8���%󨣻_}�A+�P�|Ck�d,�h�����z[��EG,au�!Ĵ�b'~�T�� .Jdl��b�o��y�6��:�w�fW��U�3�Z��q�����h�>X�>.X?p펢�`��jYj@���2r���x�}%�	F�"-�ht����Mm�|��͢�{K�q0/�g��h���2\�;jz�/�>pk�k�A�q"���}�h��c�Y(7���[=T��v��#��'7��6y�t�QGy�Mm�z?P�V������LݳU4�`^
 yp�.tyc�|��~�$�x���+ٙYߓ!�Sp53�"�<�Z�E����w����h�K;%���k�6���!,#�^I[��pXu�=o��`���9
g�Kٵ�o��0�2���|��g�F{���S40���l_��|r�?X�[ܴ>�s�V��>
�ϥje����j#�s%�h�A�l4��,�����C��-���):��醌~p=��0�m[鶫��n�}���<�����J��7�/�i�P�Mw������p����ڋY��]s]X7g���
h�ǭD9w�����b�|�0�'�簥���ˀ��>��+��.����P
����n0r����2��~,9�U��9^�RZ7j����.��|����l��	��Q+��d1ҾW@}oA�#�#��P"FM`��զ�D����2u9������Q���O?�]k�U�/�Q�ibqz)ٿ�#:�/`�\��������}Bn���'�v�:����>�u�e-�5W�J꺚�#�E��4���w���ڊ�ZyJ�-���L�X����V�F!�����"Z> ��01�j�8�rNP&��N�҉�w���tU	3q�;�D-&ݼXk�9nu���J����r�_tn����
O���Ќݽ\g��"'ܪU������֎WliU�nD}���_vx���],�i��t��]�=�$�<��/�&��S��r���*8*
��_!���A�3�q��fP�����U@Ff�:��C�a�04"e�d��\Y�γ$c��P����)�T��q<��o�A��),i�{9�p��~e�� %�k�f^��K%�D�u�Y��ss�HB��2���YT�m�����--��2TI1�w����J�!�N:�5�����0�	�p�qv�P���g��"����ƅ���L�{1�fϯ�s5�)BCU��~���4�s c�B�!��o�ޏ.6�~���|�o�SK�&3��,)���	GYG�� ٤�Te�r�׸��Fa�'g���:�;��b-Me�l%�w���&�m����"T��:�$,S?e+�
/�����Z/[�:]�0+M��W��M�ohH��L�t�fw�1�H)D�j�b*d<$�	�װ�r�N9�h�O����yK�y}sʋ�t�� �7�i���-׎�d�>DQ?8�g�l�����1[#f��M���2����0�~���7��\�;�p��ʱ|��?*��#�̕�?�D��>�T�O��{�� U�3M�>=X�$	T[4
��z�����9-\��&���$�d�r��8 rrH�{�'�%=U~�C��9�VMc�+�Џ�� ��q�g�F><�h�*�q�l�+�D7[�V��g�Q<�>'�H/I+pN�OOYX�w8���P-ZZ1e�,�F��t_���9lN�����B��� ��\�!����4��c���K�G.�י�����N{���%��o�FǙ>��}�x��EvM��N]{���g��xA������x��N0����� �N���V�c<�,.����s��(t
2|[ṣvd� ό�l�" �S��ڊ�#r#J.FPnە�BoZ����T'H�(�Z�I�3��8V5K'C�k6&�?�f�g���QMs�F���H���s�?�h�s��%t/#�*$[�b�/�^��yf�>�c�R�L��=�������T�[������Ȓ���F�#KF2G"�v���K�2*z�gj�����I.�῾�Ks$;��`Q&�R���,�g�Dʙ�#�����:�,J���>���?�`vD��c،UP�$�*v��ܨ�C��K$tprs\�Q/�f��u0Ҩ��[����Շ�����˥��������S�c�.�F%��DF��3�ڮ"̶��EQ���T{H�
*t����~ǹE��}	��\�Ү�>���_)1�LD��P2���ڹhDVQ�[~)D�|����T�49븤�R�j�A���J��^z��@��ׄ"3��,�8��d��>�坍��/2��Bě���	;�%"t:}��I*	�`�{�������=W�)ȽT�����z���2><Q$��<�!�iSF��T��ڝH������B��Y ~�UY1���k�G���*��z��˓�M��-t�� �os`��1pYI�$N�̫��Ա��{�v֤b��,��C��:�T�pQU����c�i�Y�h�Z��#�$UC�}ٽ�bU�K_Q��d�~��v�s|���Q:���C��[����{5���FxٱD6ʃk�v;$\:���yx�>렉�����8���zF��N�C��W.Y{.�t�0C!�j`�
�.t�ie)�U�tڮ���_D()8Cʰ�ǵ- p<|��Ƴ��;��}������ͅ��s��3q�;���R���"*v�
���G�P�c}��P�.t��H��Ʈ��p�(��-E���0� �]�]����ǁ�4�@��[�y�.�a	paO�n=f$�C�c�.%�dPF�a!�9s�ǣZ��	{���t��5b�9t#�{u�J��@�<ǔ�z�־�܏~� ���k���y��F�Aպop�%
{��~%���C�^���A������ԅ�J��7��gl��9�i�{��������N�ԻY��g����297俗 ������e�������?n�n��-i�x��s��>f�òuI4[����F�]��I��|�x��G��<�H� ���%I�<��i7��	O���D�*����W��H��Fv�����>mwF��2��̼,�I���|�S݉t�X^j�aG98d�I}r�P���nD�}����W�N�)��
�;Ưm<�u�wԆ5ۙtЗnCK��s�*Dgj� M��~/Ţ
���*�sYg����j\M�	�{�a��~`����X�[��o�ۘD�/y�2
�[_Ę{����'�mS��M�L