XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����
ݸ��*�ؾ5�K��/�G���yL"���7�Lנ� ,�b:n�mT���򣠧*��lR��npU�=���� �i>8���w@w)��q�Q����u�ǡ����LfP�ގ�J&H���&��஻2h��7�t�ԆFYL�}��Eʗ�*��Pa'#G��dK.�Ȃ�x�'0� ��7�����.�'�6O��@�M݌�[&3`Ƌ��{5�x�]�j;u��4�f��d�����[�¿o:����za|���uX��ܸ+n�G���|����!��� �����\���;�����2�6�~��8M#�k�/�}�m�Dp�P�A��˻ˏ��l�ӎ���s煮\���'k�d�؎tm9��� N���0��pT�0<i����l�����i���ȁڜ\�wɐ���BmZHY�7��+��jN�Z����-���d2��&G.��b6F�뀥�ш|0�S�Z$0ƕEţ6�I�?/�sùy�TH��֞ '��&|S�y��|˧��{�9`�z��n�Cxϻz��LO�"@6� ��'|��8��z� �i�"	�ӕ����F�%\ �|������Q��ڤ"S$
������6�y�74�LO��������]�* �2?DL���o�	�|�rttМ���������j9F���o(iͱ��3��E��=<>�h����/<��W���r�Q��7�P6���V��a���4�
�iq��TN�Ur~�S�X$����k��zޟ�"N1�wXlxVHYEB    fa00    2a40h� ������V�9�k
�y�ܝ�[��O��z�!�?Dm@U&9cI�{Z��@1W@��[v����+m��	�W͵i��x��������P��\E���3� (�gc�O�� 2��D���ݠ��N��T}�$�����ˁu1Ƣ�܌��ŀ�l��Ԝu)I�M�=x��D��C�Xs�$��g��X��2��}v��>�k[b����|�v�P��:Z��s	���7>N(�9��Ǿ�7��X��-�q���E�R�?������L�KG w��
��&(���=t�`q�8nt�hQ* �r�5��/��y]���O_n`Nu�.^����S�?��ZM����B����A��q��k3J�N�P-Ԇ]��c�9qFT�g��^�@L���Y���A��9ߞL:$Y|c>	��xѵ�|�a�����:8�L5��.d�v�ζt�b����^L�
\�9��R�� l�kWX8�R]+�d,�~��WYxx}Ms��u͌NQJP�yE1�J�fo�QƐ};����p�Q��������ִ��'Z'�%��ޣS��T0g$}s6E#p�I��@�ݢ�o�̤��� ͅ�!i2�z�.o����V��C�=���>��������T�H�7
��m˻4z�D\H�$�~�����637��{h|.���f�:f�6%H�]�����
�١������`>g@�˯ƻ�j������k�A��u� �\h /W>�Z�
�(��{������J�z��Vn۔?����>��n�G�Q���#���hYP�}�o�������G�`B.��	��׫�����]bU���Z��J�^�@F�#B|�8�\�e1R��D
����L�:�NcP����o����A���D.x��G'�@w{�t!b�V��U𫰫h����wp����\�7� K���6u��/SA��Sc!䘜Ҍ�����-��M/W;4��O�rR>$�Cw�:�LW��U��E##�0{3#��hy���z)������}ͥ9�qV�f��K��t�:P���`_����P�{@�͹?!s�6lL�CҡdӐ a@g{�}
\~V�j,U+̓^�7�o��6��{��^ �9&���"�	��X}�U00�]&N~�����pډ�ELXK����a-�p?��E��m\P�m�dz���-/���߶�f ��UQw��YN4�e��w#J~3f)�*�����I ��ֳ������ݭw?xgf�F���N�^�c?���h�6��&�sv6b��e1/��!z��\q;�� [�c��+�j�	z�ld{r���[�}L��=DU^���zY
:(�d�df"0�~��u�3ь2����u˙g�d����bv�m���v-�UCV�p�6�7Cl^�9"ƴE'2�f�d�J��A_�h%����^'�=8Q�����9P)�O7|eϰC3Ĺ�.��i	u��C�ş�$�н@ݭٮ+4�O��Tѯ�8*%���&yAӮ�r��E��d����������.#r�ySR2��̵���Zo<��^�������̨w��dx�f��i������>P�l�7i�6rtplsA6.~?�)�C	z@(2�{�����!Z�qI	^��2�(C����j�lE�ى�u���*�
�
�oki�Qb��½����	������S�N Pr~���zL�K?Y������J��Z?O�90b���AXJ��"�����-�зb���rp�!���c;SMC�Y����v��PʡǗ�z��膣[����c�����Νg����Z
\���y � ����S�r;�0�lH`J^�}�,��R.�ck��~D�#3~��{ފ�
l�=�R�����^�e�T)#;�`�$�A�L��I��F<-���P�l&M�|�h����Ѩ����r\�����&4Qb"�Ws�7dL&s�T���.ԎI���X�+�`���8=5D����G)���6B��8v���J'���K#B~+�>�a�	�*]����9j�����Z lܹ����(��G07X��_�70m��Z
�ٱ~�;�����U�['��QM/�6{��8���d�����N���s�ֳ���wh�8���!/Am�)s�%�PC1�W�l����@���챬���Z���b�9������A��r�y���'WP�	*5�Nw$hOHvE����3��=&�%���6�w-u7F����/A�
 ɷ�>�햹�i���+�p�Zٗ�a�c S��J���h���-ˑn�:;�0p'w�^�`]���b�ya�<	����7��T۠�ˉ�Bar�I�kNٳ�y�:,��b*!9XS�M,M�u��&0��>�����x)I������FI��x���]^���P�i��~�;"���|�F�1`�����!'�e>���4)��%�9GZt_ �M��h�I8�p��=yjQ{|��=��+�����b�~5"�m(�������£!J�`Iwl�ç���u���[δ�������!�ep���}�n��������"�ރ�!�V���65e��	<iG�����t({�5J�&��7�Un��U��i(�����V�,��Ia�r�I�d���Q(�3�3���y�񡧩o�u���U%�:��~1v׬�%2zw>��Le��kTu��DJ��x�oǎ_|gWES[O�Rl=ۤ�9��9L%J�tQ�C�4��'�*�.���D���E��=֭�gJ����]͊\�c?� ��o�{G��k�Zjw5!g�<W�Q�d>Zv���g�z���5WJJ������꥓��8���:Ӧ��VDgudw�˾���I;�į�:ڽ\��b��"�����5T+FH��&uԛ�e�ŧ�:������oӇj�����y�N�7�'����"�l�ҍ�8�!�]*�.v��^�s"�ő1����ƞWǑ�6F�*TS�3�S][&���3k��K�n��U��QzdU��P�W�hP>2���?���j��t�:�4����C�R�a�Ͻ�%j(wv����!i�Q�z��<cVI���c&s�G�����!
��udJ-�b[K�2�ұr�Z���(�N5l�WOXq k�@�(��7��_��>+Is�ܼ+��70M%�3�'�T( %+F�k�kl�B��u��_y����Lj�;��t[���N�4#��G��_i,�{h<��
*�X�Nv�����T��Y�T�iS�S����^K+]�7�h�۲7�Y+X��Z(!F�TNF�����D�ɣin�L ���a2���;1l��2K(�=������u�l��B�M�J��dnȘ��؄9@���q.tf��}��_����%�_�h��Lf	����C
 5%`���F䚚)*n [�T7��ߩ5�꺹"��a���q���9�\dzQ��J��Qǭig"�lqϮ���4$C����9�������"U���Wa��Ͽ�D�P���})�&�)����������F�w�l�-����}do�����]�
�=�6t�+VӉUc�3��N0`��NH�(�(����X�ޒoU4�|2[n��nP��I���+qcu�eAղ�� a,̯7��h��H��Z���'�)�i��24G���{�I�mR��x�|Y���aio4��ʗ"�%t���r� �]�f<������!A��Ճ8WG5�l���rX�X���8�1X�%Py5T�xtZ������4%��W'���F?�nu6d��OB��k���1JQ�^�<��R����_��`�Iⷼ��!�%T�v@����aO���?4��������B�0����t��t��B�^:����+P�ū�*:b��ı:����h\Xq�4��\�!�ϸ��o�s_��A���d�m���7Xy��YQ����"��q��JeB��q%�H��c[8-q�?p1a�^�o�D̕���!>VH�A<�2�����`�O���i8K4���'�7�a�e�������f���1�@�s_�T�h����8�Ʃ/%��xB�VY���!OBH�%1I/�<�ܤ� ���Ǻ	RPɎ`�Ҿ��B�8T�� �]�'�-��iI�h�&�C
�N�	�"W�$~�;Ք3'G�B�Tu�V!�`m^�S�-cv�	����(v5u�b���	�kU`�Ys/�޿C6� *�^
T)X�<@�vF>�xOX�Lx�D�S��7g8L��EYt��6�����dd���������+�� xa�_Ob��?|ܓ�$�iR�Q�\A�k�0��u~�S��I�O���r�m^U�o5�X�Nc\�|
q��E���g�s�Fɑ����X��ǟ8fFo�XX��YD�;P�}"�<��}P�sK���B*��w.3`�-)S5�;��Љ�DPI���a�k��|�1r|�� �W�����"�kT�5_�(�(6XcL�6ٟ�S���x�WQ~	4�|�Ȍ�k�8le�K=��`����K�����)��k#U����,v�0R2����xf>�˦Ca�N����)�H�ـ�����#�X�1�܋OŶ�٥�<�h�3dR*4��;5y-���/J��b�7�R�\1�/c�O��^l�>|V�}n|�>�d
�r������ԙ}���{�B���ڴ��q�W�\��2tb_�Q�t�J.u=���!��bCA��^�$����s�Io)�4r+���Qa*��Ρqd�z�}�p�/؉��u-�gqg>���[�O�N
� �h����)(E�8a2��/�:�^�o�LtY�?=�m1ڪTqI3���1yg�R.m��B��=��|�(]���p(�g)�$�'%G�˵C�e���gi�J��4�y���=�{M�#*I�믽P�L���a�<-*-=,i﹟�������=P����:�^�v��N\�Hb�'����_�)�R!⸳�K����<)���DrP|s%�j#�����q�T}�H_�-U�ԙ�N��R��X�\߅z@���m��Bw&
��wBl�rJ��I�d�*Xeؼ��~�A2�c|�[r]3t�An1�
�?��ǫd8�l�z�x�(���� ��j�v��;s�;���s�s����*x��YI��G�8���(ϱ�ꠋ��W\��JKB�c��r����EW�ae��Q����\����4%���F*-t�Yl�ɜ�h�@��f-B��gq#�Y��Ĭ���ɵ�xf��������.�9CT���5���U�ë%Z����n�/aVd{��n0'0�2�j�q����]�}���b��=1eN#�%7��E�*O�w�VU ��}��N�v�I��Q	�~ZbNi"_�����l9d�41u��T�tS�W�����2�'[3�A�"3�D� �����o@B����P���t���p�gO!� ��t�Ӈ/�#��s@(���	�Mc�ͅj�5�"�b�f���"n�9���7S��pi���~���1�t�&���v]��fb�ω����ݏ@�z I�O�3�O{&�90
��z��s���/��ok�<��wk����`����L�a�>��:�1t�f�c��͟�����^�京M�*˰�������y����T�	PA�������������M���a&࡛�E�=��ՐQc�ll1{��Mt��7Nފw��)/FH�I2ĉ�`���� ��,_��:O��}t_*d�lP���B�O��������t�Δ��Y�0�'Xif5W#~�띝t�6�ߘ��8&w&���6���|D�Z��Z79�qhrh} >"�����w������Ӈ�[���:��x��iQ���$@K���|D!`f�llR���a�{6=�v��
�	ų$mr[�TҸs���`��L)�~GBR=<q����1�����4���安�DU��m��=��� 	B��-�ڔ�C�e!�ҫ�1W�Xa�qP�J��z��[�����@��Ʊ�Xs��)���	�g_�l zW��&�C#	� �~G�$�mL�mB^嵲�Մ�0zG�ffG��p�]�.}Ԥk:I`
�&LI�����<J0�;r׸���[=�*f9���9�A�=�y��,o�t�ȟ�X����bI8���ڭ��*�?�E#�R�*�؋�.R9���K�̢wpgz[kI�����r����At�B��$�Ծ����n�� �ҹ
��]Wv�^ ��! �|�,|�	�D�{�����2k����uK�*g��0XeO*��*�?����hp�S$��_U��3����MG���Z9��p*M�z�Q�ZН�
��0�bz! ����޵���H=��:��G�]�ڄ���h��g��ˤ�?���6���f'�1��pVp���H�&T|F/�(��
q���guW%�W$���� �6pw��\T��䨒x�?���By@9\���&>\�b�ӏ����~���-ꑨ).��#��K�n��Qڌ0T���6(�R�㬦R�q%�u��b_E!z_��[�+�̯RW����s��� �xD�M�+L��ۆ˾3��ۄ�ٞ#K�����B��9��H�F�o
�X(<�	�R�]�)}���m�3�پ����/�;^E`k'�^4����)mKV�����xUbÜ�T"���א����Җ8����B$��x�w�4������1Y/S��ڗU̠�E�U�]͗9>���l�Q~i��-�Aer��!lai���
WF9�И_�}E��'Q��U��Ԇ^�X���d�
����������.<�,y%A����DR1���J���6�`r��IE}��qL�:β����c>�V�zG��1�
ݠA~ݾ��k1�QmHc;������ƣW=
k��kE�ͬ���?F�0s�
~�9��_G�`+s�檳ߏ�Fv����Jl�M����d�i0#���
:��$�[� ���cZ�y�QH9t-Bm��a���7{I��8��Z% �C5����Y�*�C�� A���Fb�v-�i)��ލ�[��u���Ѝ'�j�/�Q�H�C-�j�{c2/�d��7S`�T蒔~�3�L�����?u��e���
�9�#jX��&$m����m8&�J�a�w9��H��L�f�H���		$�����Hf<��)t.�d�b"�j���/-A~���s�Z��qy+�w� *rn~�i튤���7����R�>9����_6υ֫��)���D�~x<}�zk8;���n�J����zQy{Cu����s޼����/=�`8�y�l��ِ�7v}�����r�&��֟�ތ�ܜFb�������+�!�G� L�t�FȰJW3��q[��t�1��6>0���ŷ�M�I�HFg���i[~��釜DLI��z�ne�ӿ�h�|�
K����Nt�,"�J��<�e��6�!�_��g6����4'�u��I�&��U��e+;�1�����������D�-?��6!cF$k�v�o<L�|O����_��j��~A�W��O	�L`+���w}A)�T�P�a�����*_!)5t�i;/e]�J�dqT�Ls�Fpm�GYv�S�i�f�|es����x����_��P�R�Y�" i$k��gU�C0�W2kFU���Z3�S�er�t
b�%}���U��I��4�Z��s$�W w���Q*ҹE&��K!*����?S�n�+7��$ 5�:� ڹⲟ�H1��'L�����I7��E���x}���֑MRu미���WK�gP$"��y{�F�'o9����E�9��N�ǹ��+B��efu�M��^�V�
֜*�r���:���v�.V��� ����լ[R�e�\G��/)>�Y@6�k0^ѼP��P����=i`#g���-�;�U@�����U�k��f1�,��9\T9s�����i��knn'�~���B#;ɏ`N\	�~D}%���9{��܂��A��G��F����"�����AR���/VjP?�V�ؽ�hB`���`6��N��hŗEJ`�0���� ����'����C��S�ꓨ�K5���e�ю�=V2r1�\�݂5��?RkDO� ��	o��J�
]A�,P�M�q�&T��}��ztBlPElZ�P%�U�����X۳v�D����D�o�������M��3W"/18�#V��X�pV��������}�d�#���?�|��s��l.Nmi��v)�"�^���˨��?:ŕ=m�D�,���4G�SjM^ ��2����Y�T�`����\�iL��"}Y��ʃ>JbVD"x�[c�xپ�5�PGr�����2]O��Z9P5]���,�ҍ�$|�u��9'��<f�!��s��.�%��5�q�=�_��q'k���R�S]�����Ƹ���<���`�C�f
�9wl�Z��O�D��!�Tk�4�/�w�^��l���B��è>߆�����Wj�U$b���q�s�n�_Y�v�)�bt}'�� `���
�
�>��_/R��#��0��ňZf=$>��"��?�$���E�.�`L-fs�.�&�*�k��&�
&y�2+��.ɛ.�^i� ��1��י�I�Y��m�b�X�3w=��<������"q��71�&i�+��qn��:n�y���-N���w��/9��]>�6���<Ցg�w���>�՛�B�PTjlF�\qXtId����.��b*R��N�KDy���5L�^A?ʢa�T/�a3SY\P��� �+{�R��-�H��E`zj.�W0t>^�3;�)��w�IN�#���.^��ү��ɓG����Ʌ��q������<A��6�X4,ơ3^�vD��m"iZW�-^�Z�k/?M)j�u:QW��Z�KF�j��Z��/0Ib,��haL0��t:��;�ڻn����cH99"��Py���D�7SF�6���H}hO�7,�Ҡ�*"�ۢ����TjK�D���ou��S�#�U��ar|�"�K�z.)ƚ���6[Y'����;�g��U������m�+�]����$� ��a����!�[YLӘ[�"�������jV9˫.f��ϖ1�$���ɏt�� �YC׾m�.3�8���|.S�b�d���o�"�m#2�z�Us�Z#�:w�H�GoK����'�q���i�Ѧ��ex�kG��RE�x�o\2��7
����å���v�`'�V	����L�Z ���j5��t��>u��;1���"g)�EI؊=�d6g\>���Aɳs�ZW���̣���oU6k�-�r�C�gU��KK�b���8��;���=Aէ��#P�V��ҋ�#�a@���OK��t�w��R�G��v��
�zm��-=�9�+I�v�2���7��296�^�L�m)'����{G�U:8�ݒ��-a:勞ǧ�ur8|��u��Y�o-:]Pұ�l<o����P�ΝG��6c��p�5���>U[��yy�`�i� ��̇u痘qO�x�؝	������A��T
�D�IDWex�-Cu��gY��$�.0|��j~Ud�M��MXU�k�u��O���Pq��=�Ҷ��0�ª�M��X6��~D�Y�IBtX{�p��v���Fs������B7�]HG��F�)W՘�Ȃ��Ӟ��f�%=� �R��BW��4me��z�_���,V�h^�: ��z���iEc1eTm���,�"����+%�q�5̟%�6��e8:IY�+���+������q��v���Q���6	`���b�,�u�(l�(�KC�bl#��(�ʠTf���\L�Y�7��@�w/��P}�!�웜@�OC2C&G��vC�_��)�k�!a�@�Ma�I��v�*<עͯ\1yx챯�=#Bpq����IO��&���9�k�w�>@��c7	 �C�ئ��l|H�RU#�Gm����.��CM��_�'�����3��Y�Q�r�{>m!�w-j�Ȳ�4�����I����rs|�t��m�j�>�J����C"�V���|@SHW�LڨV�\߉ٌ���n��?�m7��E�yew�=ka����o%�S˔ގӎ��#�u��.��PA|/�tſm&�i!��InL9�~�V/��~n)=��~�$�P��E���_r��T������A6�<o��^Um�O7ѡbY}z�k�ء�I
�(�U�D������1^d�Q�r%p6O����C�uw�B����ǈ36=!")-��0��}��B[1H��@"��e�Z�j �徜'&Dސ*�\�\$�aL�v�*�&ڒ�jy�x�4�삲����`� ��l���P��E/s���=�Y^.�_��P��*��y�+��-N4[F���|�4���+?z%�/!m�&^�������P,�y�n*xE;�:� v����Ǘ�������1�Z��\ Jx9]�kT�r���G��l�Ԑ)���b3��Pb�i��y쀡=7e��&SQ�RM pY��޺H9�
�TF���m���1b��W0"S&u8�١��rժ�b�<��ȳN�|?��UWK��h�(�D�<�eZ�`��I@��L����
��DL��I�*[�������i�:q/����H�l�o�	/�ְ�^��L�]������ͻ_��'�v�Mc�g��ތ�嬠��s���k|�c�-�b�C}��r��Gw���b�f�+����B�,��M_2B�G!�XlxVHYEB    fa00     8e0�7$j`+�IۺĽxV4�~�'��K��9
jh���#z�����͞��T���Vj���u��;>����ׅ�T�쏢!�	�z�����j1�An����0doj��*N���@!�,lݫ�G��g��e��Ժsx��vg��[��	*�0y��1�x.0��D���TN��A�-���	%��j�3��m's���.j�F�E�şoa��RHދ9ٿ<�n���ʀ�	g��Fׄ�iP�%Y%>-�>��b�ה�|��v~�u��ܡ,s�n�����9#��3^�aTh�p�aV^��D�L�B���_F���̒.)
)���R�`���o)�F�>�����ΐ2A�t��ɋ��x�ԙm�y��
daƹ���~�����o�Hjr�r�f]Ei|�N���B�z�5q�'�\V!O��C��MRې��S��j����S�l%����{@��m!P�|��GD�h�/�����ŊA��=�7��w���:��@���e�U~Q��Ԡ�a^:�vuJ�PCxz�/k%�l�r��ԫ������*�1�����7�9C�����j}�]x���c���gSA�LˡQ�x��̧י�4�Y�'�$~�V��Q?&9�8X�+���'�($gC|�7Q)�ˋ��rR�Ώ��7�1�����k���(��$�5�a ڨ��%��V!x��3_d�p2�0b�� ����p�-c�E#/�-�(��#1�S�!���mʼ��<$�Ca���klm Ab������4E��R�Cٯ�$��] /04�-m-�Z3u��������4��F�J��3(s�X�¸dM��$j�|��-�3���p�f@̄R��r��R{0�f�Fm�gE��V�V��g{�����i�		���u6�+��������*�o�!� �уx~�L����a���5�zzkf`8k��ܙ�f���D�ou(�B�0r
��1� �}Lf@�-�s�جFG��o�-C��ݱ��w�e�r�ꚽʁ*ӌ.�&63j���� VH�
���֮��F�ܤ�Z�:����O�f�f�&G���7\p[A�l�?���A���e�5�zd���&_�Gvų���`�����R��_G�Ir�k��J����+�Ês�p�#�o�)��)����བ�Z������\��Q��1\�Re=��0���-�L}�7��(�Q$^9s�A�V�"/8�/��o{'�H���L���J&�|Q*�/�?��L>�,��W��^2tW�{�ԗ��GV�Ns#��ўQ2*,"�HR�|n�i���2l��bm���H�Z���!��_!� 5�%@̚���G�'�ꖧx�vЇ��M�U���`�KTE�/b�$�� {։������a�x�<�@*}#G�;ha��v�W�(z�U?>�3�F7i�e������Ӽ���z{�X׋3=Ei�a��DP�fӆ��H���r�ĭz�;�������i�<�9�>�����ÈA�FkzO����t��������ԮO�^^2��}y��������qD��J��v�P_.|o���( s�8Y$��pÖ��
��R��B�j��N���r�zL�����X��� U�ߝN^[�y��w�}�M~�"����A��b�Y�2�?Tm*b��/6�/m��ϟb�c�0�4�UD�����E�0f��4:�4��pG�����4ѯAj��L��l���O�_����M����\_L����?6���X����n Ԍ�NΨ%�4{a�X���^����Ij�2�����������|A[����>&���G�g���ƚ�N
�Q���)vŐ�`��	����t�h��A��-�Lf�bǠ"�	k����e��@�X_������:�k�S�C�f������
��ƀ�v�+��`R#;t���,�l8�^0�S�yc)�ǪZ'B�p�������g�ݚ3�x]�JIHj��J��I�/���Eﴌlc�'�L�ah�l�Q�aaCj �ǘ�`8m�;y�4�����5ԅ���=Ɛ�S����9 �	�k���4�	m�����a�W��? ד}�@�R�4��F�5qkV|��4���j��r��jEz>�Rv�z��C/���|4�$?��1�H����S���k$E@�A�->���l,seZ:VS_>C}�Jb��}�<?Db�P�P��Χ��$6bW���W�5K2��!���&y��=��w{&���:XlxVHYEB    fa00    1110�R��o��m��Ӫ�����^@���L���ȩ�ZN9�5���k���)��ͯ��\�zeq�Ĩ3-�,a�����o���Lk�w'��]M����}>�M�gaă��[���KDg�i9�����m����(.��i'�-�]S^�9C[@�e.���iW��;�JQP��q53�Î�{V�5��S%>�����D%��|��f��m)�M	�c�B=�Cƚ7k�ݰdVX�P)6yp0��	ƀ^���_����Z��O�P�'�<`D)&��"G�&�:�o�'t��ӎv��������(2�'>.]�o�㖘�d�A2.�󲛵b���O�vx�8@2dz��;g���?a>�*ˠj0w�j�>�Z�?CH9ĵ"─oc�	�v����\a&��&��E��Kc�K��a�׵�dp\�b5n=o��l��X����T:F*�QJ�Ciwr5������>����$~]�"�.���\3��z�O'ك����J�������E����|���5�K�+$s�˪�7���!���<4oC�;&�D�K�:O�Xt�*Ո��Gw{��q�tj��h?)��B����y@���D��,�(M&>S2�᎔��W-{���u��~��"lg��W�M���nG��?�xP�4�8�s���%�빐�-���|FH���FM�����m��=D����$�j�zX����C*����b:�=T&r:Czt����(_�̉��S�b�m���_��I���M���!�8��i;kF���u7,@!�S���+;�^�z�e�S�^ݚ3eR�9��+;(����C@� gTfµ�6�b����-}`����	���x՛fsU-�K�͟N�ms"?i�/�?ӫ�Ǳ�#����5����HQ�v��]�C7�敳�l���g�)�m���a�%\�A���-)Bj���$��7"�>��Юpo����g]�գ���a-�tE%��a.��y^Q�\�h���n��R�(׉6�~dJ��:)Z��.)@v ��U�02��H	=��G���~u����^&/(������4�bL�%VX�RA
EF���(j8ᰕPJ)gc��Is��w����i��@!B��� �����$���Z�Ґ�jl�	�.}��=:�ZW3 /��hl��RF�c���	����+Y�J L	��nXm�i�&u��Tƒ��)P�}E	s.3�G�m�S�2���yl�6�<��0h��"]^���]g��sN#<��z9(Li���B��3b0oY��۝>���6�~b<��uE�(��c9Z���!7m9윛�4J�*�z�2����i}<�H�4Hr�0�߀�~���KѢ,,�ʪ���P�p��җb���>�QL|�R����B/�&b��^8�v�>Z�1��GG2s����M_lP���2������wم��λ1e�=S�a�G��/+�jo�0W�ޔ�;���N|���V(
�4$*#@L�#�^X'�����c�vP$ː�N'���`�������4����$jr����W~�Ƚ���+�u!��k܈�A׹
��?V@�ڶ�9�C9�y òXFr1������_*4��b��pNQN�������yr�h�e��+��7|�Kۀ�PL�4�f8�y"�gS�x��dZ:�X Z�9d �����f��ۛ��}�����<�-�'&���9��K��-��A�^��Z��=Ө���7 ��M���r��L�"�LH����[� %  Hs0��|�J�k/˰�B�3.9����=����i����	�M��w_��@E1E�۸KCBs����t���*P-/1��䍬�J(w��+U�awr�)^����˷��j�>�9\'��Rf#H_�#��4�N�]M�b~� tt\�>D�j�S_����3St��3�<��}!��j�D���Eh[L=
-��$\R�+��Ӌ���OZ�D6Yq�ϑυ�㳊�A,(���׏���gg�������T��.?
;�ߘT՗@ 4E�Ǚ�b3V�O�?�?��G+��ź�V񻰂��cEC�s-�J�RRm��P�v1��dI�k�^�G��`���1E���Lq�=��D�?�٣��}]�&��]�҂����W�3��ח�1W�e�B 0�34�_껍�S�,i�p���6�ur�9��
�q} P�璹蘥�c�B�y$ӤG��^��*M���_r�1L�Ii�=�D\�O��N���L�a%o�̚:��!2��h�"q�p�X/�%mD��q���c^c�{���Ⴣ�?T0?�ʗ�`��n�{��a|���ᶟ�����e�\���WGZW-I��@�E.mU����յ�e����T?�=9��m7�^֍��URï�c����mvG�_G���0����щ�c�/��c���jȭ\S��s�Y���(���k#�9�V������WU�5��A翂�֗�Q�(]K��k&)QQ���k�w�a��
���Tv���A�^Ɂ{��O�{��e�"�3�W�hk�H?�M�(�W�L�~t���։ Ȇb�o���eYZ�k�BK���Y/�$��U�T�1�d����:�	[�W����l�[��Ŋ`��X!R����hm�3�,���0f4�9<�U�0��:+'���i#���t6�d@lYo��W�D�m��V�F�H5V�x�4V>��6/鳎�9i�U��bG���R���-��m,j�7瑥�:טN��oi�$�ب�АB<�Q��jr�J��"pr�������Ej�\����]��2�0!tC�frҥ���*Ph�����86� M���L��=�Qxv*�%y��F���G���P�+���
!)��_��!uo^��6��R�������U�r�ph�|r
%tú�K@X�.6^���^���$�F�G����F��	1�����ώ�G"`���0�M	ݺ�H���=o���]x�e*J��iG:��f��'OĬ�+�O,)9p}�8��%����N��x��j��� �;"$�igz�q���Tb��4�DW�/2ӪJ�,F�qA�";nvo���O�L��b�f�a�/��|��?)(	󥰒x���B�శ��:!��'RN 0z��T���O.�8Q��C�;�]�Hd�{Y�HGbl0�-����8&�Ye�/��\���E����Hc�c�-Iz�?��^X�G�Xt���Ӊ�t��M���w wVu�I�v�y7�5Fe�r�$n���J�T*��0L�������!���Ux�zt�5Q0t&�.ܥ�o�!b������B�%�dev�7�����>�������X8����b�V}��:H�����(�`\�5}��}L���u D�Þ ?��a��<f߿���ձ��Y�e;�O'D�SC�{�$��u�,��YYl�Ch�/�qDk�@�M	�g�c��9Z���ĹK*��E|�w|e��������k�_�KD� ����<�Tʥ8��t��������$��L�ف֢e�iKɝ�����m!c�ݒD�Z
�G`�Xq��O�_S��x*�t�m����;��%;�Uj��F�v`Œh�fX�$�4��7A��3+Af�E��vR1e���ɬ�
�ՑPJ��(IL�ܲ��O[�mb��e�8��VF'�JR=�)�5T�Źe7�^}2��r'=�f笷J�:������X:�[fۧ� q3������5&2���2��!� 2Zc�ck,㎛�8�#��s��j`7���	ַ�5��砈�*�d��qӓ-;�ғ�@ݙ���_T�'A�0�G��Z�G�,���O0�0J�m��K<��u��鶄p� �)��F��Q��'N�G9��ڇ��e��얺��s�����dE>���Y.�@!�k�'�j��4�=c��!vL�";�j����K��2�\�^��],�U�58D��n��7�bP�@Y�YSV�]w�Wlcל7�cQ�*�2 �G�V������}�qt�Щc�g�������Q�4!v��0��߽�I�ǽs��O숔�ꤎQ_�H�"!�+J�0ɍ�GD>��%4�o��w�mC�1�9epPi�x�q�D��0]�}��b���L�!���	�.�T�9y��WW�`Yy�M��M�P*�{lwKcαQ�_`Q�%s@w���*�4x�83��3�Ĺd�����m��caNK��Q�1���LwI�F��m_N)w��pRjV�8�χ�0�� lb��#���j�U2��V:�-�]����׌'X-{RLtIk'
����%n�׎a:�\e
H�XlxVHYEB    fa00     ca0�JUb<T�0��M�]����".���Kkr��o�q�s<�ف����HK/KN�%TX����k�'n�+�x��g]V�(tݠ���t������i��8UE�N �h�JL������e��	Pٞ	��z�Z�\p:e0E�y�H9��A.έ�z��c�%cb<��i��Ùvi����vA���S�WF8
9')����`��e���v�z����F�iUIM�g7!�5U�!9n���nnTYIcŋ�(_�t�V�G6�7���������EQ�tg*S���4J٪��bȾT�Y����+.?w��ZMuW�%��C�3R�v�L�Y`�� �!q��}�e&��Vd��2��U?�[kp3�ʰ�e����-��Q����!P�܈C-'�W1M2s�`�;*���a����D9�W̊o����nۯ�wL`�fhA�1$�X���2�,ZR�	_�T>��| �w����=�*���;��Q�J*׿}�x�����%�2�덤g��A^�n+���|G��99yH��+P��/�m��ꔥ�Ds�l�xȤŸ�=V��
�I#�{���"!���W���
1n��=�/�Q��pQ�}�[��rR�V@|�)�2O:�d`~�� ��i[��[��M�t��u�u\�C�~�_�s~N�MV��~����vIT�A�t��f�U��D�]��Z��3ʣ�7�LV�{p2���F����-������yP�$�B���im4O�{�?G�{��2i8g�c ��Yg�io������v:��̈́�	�\�׿��\��/F\l��0���ܣz")R���$�!(��� �v�2h��Զ�G2��Us�{T����q��
��8��9L���0���Yܶ6S?)思�:O���!����)���d��'
26HRw�tf�*p��z���
�N�M�A�;F�2��l��&*��<Ov��Y��Wgq�]uw��Q�������^p���/Ͳ��1�'���E�	�Y�{�=��k�z݊��]���~�0�$g$ne�}��{j�^��︠0��yн`0Y�+	�M�84��Ϩ����g����FL�.6����̪V)5p)��������tx��>��2B>a���I	���
�k]�&9xyT�V�(�� �DRx�?���YK�}2s��h�;>��6r�젮Z;�����/��8���Ec7ys}�M�v�]����;h�}�_�OD�#�t���S��|�Ǖ�B�������Ջ.^,x��{hXb�����Lp��^=C��TSPmF���,{�D&�qG��];�Z�.a �D6)�RJ���A�D���J**�<�$�	&K+b� �D������bֶf���)'�1�8��bR\�1��e�pLVӢ5l���1�g�����I�$]���y~b��a���:���rS��� 
ٮGtH��\/�	��1�q����[���d����i��M���W�M�:�=r��ga4^�J~b����R��u�h�}��0�(����cx�\�$��W�on
���:;xU.?ҕ�����e�#Q��*i+�)N߀��#Fԁ���b�伩ʠ�t� my�?������xQ"�Z
P����6�LP�ox�5I�F�-a(r�7j9T�|����~��W��K��<�	��4�+� �Բ��v�S� n�4"`���T�5���d�RC���')������"�I��':�!�8Gz���Y��"�PU�s[?GJY�L%5c�8��w샶4��x�L�.� �b���Q���9�n��c*�4�s?�R�
M}�۶%���eaQ��)8h$sy��4��I2k�F٪�a0|�m�����HǛܝ��u�׭����͘%����H���f���1��{<[���/���q�U-s��Jvcտb�?���U�O���h�C����XH�sZ �RR4%q�26A�F�N�	$e�S��+�%٬�/_�R�}!T�~㇀1$��أ�)*o�8���Pf5�M�m=��Y٧G��KN��O@� ��L:ُ3c[�����h�p���H�b)�3
��X4t��iR�!ۈa*y{"�BV),P\q�}T3�H�SJJ{?����Zi60ZU
�;A�	���7���x)�j3%_�����sC$�;l>�}���|��9ŉ��D��J�TA۳F���4��� �E��V|6bF���.ZH$��ofK��=�,5m����j��"�y�tȬ`�J��� j9��"�c���j;OŴ-�0K#�_ǎ��L��'��oAy���snI3��o}Xah6uݭ�0()�]�<��';>��pk��n%G�ʚRw��u�`��pn���5�Ʒ\�I�+��"`Iq��
<�ߋ}my5̞��U$kR��\#������O{rۉ��y�-�ׇ%�D
b�G��R�)3��RC@0���w�N���#}3�����ŰC�I�A�W�_���,�����b���ị4N�g6��͸�R.ăj+�O��8��[��lf��C��s�DDמXE���Ti�,B:P"6�,�E�e�?�t/F����vr+f�D����<�5����cO��86�^�yňV*xp�� P+�\SZ��uL��&&��,�Q�=��j)<.��8����B�L�V���~"��%V]�)�>_c���Y�/��h��8o^�r���pX����#���̪]%;f�V��v�z�%AC���cG�L�V$��()���xd�`��\�妦e9道�F&	�PM߷�ރ�zǛ��iKqB��A�S�����|L�l;B-�I���H��[r�>���T��j$�e3U���-�SRC>"�[�a{ۋ����p�|Q̧��D��ӳ{a�Z?�<r�[4�V��2�'�G՝^�*!��Bw$f$X84Je�ڒ�~8؂�h
܋/JX�6���݆4\ gDK?��H���>i���b�r}�eW��ءu0�i{�<�����A�R/�:���~����䌎R����&�d��(�� �Ne�Q� t�+Z�
��-;�[Y_%q:dR
ws_N��L���>4��3VӸ���)���O~a��1u"��O/cy�r�3QЏ�	�```��V8N4�T~0�E�NƆ�+*	�&xMč�$0H Nl��8�'����&MP�<1$I�XlxVHYEB    fa00     3f0U��߽�ᢃ�d?cg�|v;�a��qoH���v�~S��p]i8�O�2��=W��m>��������Vd��+~U�R�T���dғbEP_3�����wX�����P*��1j�v*μi��sc�b�Rwhɗ���v�\.hE����cݙY�C��ٽ�U UZ�IAd�w��>��5e
a��#ly=�`[䤆+�� ��+@��v���]�ԯ[�6�`���Y�}�f�峫SI��-��,��d����b�uP�8�3�2�v\8���������y��`��"��pE�C���<���ܳLg��%��5�����o���!u��#�,8��-b��۫%���y�����p��8��d�ٹ
���j��L�#��*��J����*��
l˃�����d������"�'Q�r��ds�"�\ٗ��rV�M�v_[x�f�n��'֣�&9�
��I�k��Tk�z5�51�=��8�'R��!.g�W����(���Y�@{$���I�Rʔ%;4x^�n�O���[U���{l
�8�Y�)�H�>cu�VL��iͭ'��S���a��֩���[� �S��l2��{�s�}��Av�;��6<����\�����>S��	Ym�L:O�������l�5�8c�g����%�"���/�)n�
��X����y�v�ȷ�]����X���W��;!�h�A�i�-�y��c�K��~V�^2��ċ�)��*T�b
�jS�锕0l���.հ�{��R ��3I0�.awL���;�x����=_�4������R-m��Q��Ѭv�I�'^7���i��N��Y�]�f4�|I ����F�( ��)<e"˕�]E�ޔ�)׬<vZ�-�:P�{�����`>@a�,T��x�A�f���&vq�bg��#b�{U�\sFU�}VXŒ7�{ ��4sc��{�/o2�w3��,;�>��?dnT4i���/.XlxVHYEB    8096     b20K��4�mT����2�f���As^/�����j�z�IJ�!��)�( ��g@�A�3H��-�8��!���*݋�,���O)d��0�\��P�Zm*ۨ'���C���@<��W�R��������k�S�d&��z�w�\��D~��hoG�@=xW�����vLQf8�w`BW���R0_����/���z0C�~hVW�:4(���v:����*��'�6���%/���1/�[B�L@�����&y����4�ޏ��a 
��|�l�g6tL���)��Ūm�Xf�Z��D\^�iQ��#������w��Y9 �0���]�ePЬ��wZ�+�����Rm�����^�=ᴻȋA��u|�cgZW�'�l�/�xғm��u���t�j^�8U@�`\ېF��s�w,l[*�,��S9�Ħ��:t���KE6|eV"C�h����;�}��S0�6v��-Y�������	��F��<�Xy	���q��:v
Ҙ\[i����^����Ӡ����ob]�iO]�ŌO1��QY��X"v�3�yT�)���;\�D��6)>�a����� \9W�W�#�|�������?w8z)��T"��O���Ȱz՟4��Tvxel:
��]y�⺦s�L��7\�����i��]���5�2ﯙ��G�,%o���'=�h�PAy��A����)�'vC�))�#qX%:H6�fv�R,ܘ�~O����!#����T11��o�}o,���k�l^v���d��jBfn���U��N���(���PB��, .�	�ًYDL���׎9�:OZ�;�ۿ����We�D���7��� ������`&�N�0��2�Ԉݣ�&��t�-
ٰuv���a��YP�A��G$��=u�į�/��/�5���-�Db�2��5�͵/�6��/Ma)=%�NKjK����F|��'CmP�h�+Ly�o6�\�:�l��.�ڔ��k�te��SJ��cj�+��8�B��^�|q�I��]�@�b���7��y��,���(4g�0��H8���GF쿃�7���?��*���yH�-c�m�³�8�W	"7Tfp�����^��Tf=n'ap��Ӗ��s?9wv��n��%��W�?ޤS���(&����<Oӆ�a1eI)<���]�ȝ?�8��h�@I/;�B�;�P%n#+B�չ�^H�[���R����5�%�l_�	�̒p\���K ��i��U���?�O߰��:⧔��c�㎷߽D�̱Y�&f
2��$
`�̗��<X�eh�N�X�2?� K+�8I�u��Ŵ;��ߞ�_i�g����\D
��B
3lv�aSfŇ�Q����l>�����y�t&����c��/>c��oEg�7F��˔t��B���}y�ӼӶ/+�]���Q���?��Н9�s�����>N�:����G�5�ך.D��`�d"�[5��yN;(π)�`�р�ke��Ӫ;���)�K�|ݡ}o�t'��C%��������؀/І�B*n���_U`���ۦWܒ���S_Q>n�eL���	yxֳ�u�e��a�m��C���w���W���@�\ ��97�z�N�4�aL���ni��mW�����<�X#Z�O�7򶣣u ׋��˪EH/�0+�AK2ܿ}��$ҙ�P��m[�wl�9���g_],4�A�������E�(Yx�x���G���ڮ���]�)�t�v� �g���_w_����D��~K�|XN!(�(Z���ۅ4�7�8�}l�E*�n �_ش_��9�#@.8μU�w^��g�D�m5oo]:&�l6Y{l��$���8-q�ÖM����(wU�S�e!-QҨ�>%Tl�gA�3�|
��a1���vD�FɠlKPa���]b�\v����EW�����-�j�=K������r�|�XYS��8D�슩��>�^5.���9��| �D���14�7���9p`�Щ�l�l�*.3�/��c� W��"��x�/Kxjx}���qT��g��l�@X�F^��n�c�mI�Jy�P���CE�%���:6�WN�0���� OIj�ے"�o}��D'�v�F/+�� uE��41�����0Ak������R@�"�CZ��u>?<\-;됄5��L0��������-���؁�_U��.C��MzC���h�%G͕@}z���P��n�di>i����#mt�
�Q|�����%v�@0!_F'5EQX�͙�j0�8�p��%&�v\��a�f����S�6�
��/Vp����J�X��tA �LÊ�� Pl��4U9M���+�zi��w��wNuH�}�����G�6s�^E�mt�\lN�9���g<����	+�_4dC��ܬN�E�_��3�C*��+<��liN9��S�ɜ?~��Q:�:��	8�U���)_�k}����1������e!*�(�Ci��.�X�]9a�(��do�&"3b�<�o��L ���䠎v]N���'�C��-��Y�/��"�Y�g��!b�ː_����K�g�o{��{?աV.A[���;f�C�e/+{��Sd��xܑ�հ�Z���6B�hX�9�\���]�ʛ�I�=Af{�`�~��-�3�9$c��Q�҉����� lC�@��`���儋kJ��tCu�����h��T8u�
��QB%����}Vy�Ac���� ɽ߬Ġ�H�a�QRީug��((�/��B�_C{��� P��7��y��r����ěQ�Y
�O�O��O�֥I!���;�I'15���'����;(U��`����]��?�~v�s�i�$x�y�}