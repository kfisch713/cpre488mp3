XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��p�db�km
+S>��W2��Q �"��-ݠ�w7l�@X� �D���+>/m\T��2$4���ah�iL�y~�����y=������z�ZAg:�J[�IQ��ܚ9�b���#"�:����k��'���'\� ���H��S���R��0g����k�F֤��ԋ�����;o�2�oph=��w��-?3j����OxW�ۮ�j��!��J�랏��d�`y��5(_��k�N/T�z.�^�>���.��T�1g�����v̦��}�e���0 �U~� �Al�Dv��ܮe[�e�l�V}��ǫ������<Ҋ'��h
_���ڹ��4Xiȗ��Y�ǣ��~�ǃ�����9�?ٟ �tP4�A��g"p��~�Om>R���گI5a�Y���_�V���w����ˆ��WpQ��_t\��Wc�n<N,��:nE��S)V�lxk��7>DD���3 �����Dr�@���_?]%F���\���>永�{�X�aP$�r-����huCod�^���� ��pL��bz)�m�d��'�2+w��AM5
���3?��}ԇˎs�VF�!w��'$�4��m�a�'-����ƞ2j��&�H�0�e^�wVD(�F�"{��t�9A�!DS�Գ���C���ݭ�°h�3:��}/�w]���`�#A�`���ݮ����˩�'��l�=l�p�
N��\���7���*ob�.�G�Ks��otYq<ٿF���
�FՁ�)�ON��u�)?s���j쐝XlxVHYEB    1421     7a0�̈́F�[�डt�S��<�ͯ����"'�L�y��蕦aX���3+����!&c�t�8��B:0������ж4:�֋�$
�����d:?�k��u���
����z{0g[R��=F �
��g������ܚ7]��?/���H�8$�S� �m槴��k�Q�~0��:�]=��\��aٙtҮ���p�$u��)W�0��*eV���������"p�g:�����ar �~�qv,`��]I�I%�eIQ/����M�>�e��p��C�A6��	ǒz�|B���]+h6�#���G���\~-�f�b}d��F�m�@3��H\��نRt���R
�u=Ql�D����d���h�y�2���-�~�>��$ox��V��� 2�)��=ġzT>�<��dm���ٗP�ƺA�GxN^i2�D���Ж�c��P��&0�L}/����zz�݈��ʚ���e��� �^dΔ�ϻ`��P�m���n#1/#!]�Q�$��)���Cx�)�+ �"���q�k�z���#��1�: ~�`�FxK�y6��vk���wc�H�Ky���ʋZ�8y����I�E~@�;H��:f,G{�{~���n��n/�*u�K�<����K ն\lI!ӵ��~T�C)r1,D�����i�+q�#J���5�<#��B
4���Z�_���*��[�
*�X�Y�S.��A�_ؕ�I��xL�q� U��rI�ơ�?��Q�e	"!���ݜ�B]��pU��&�˚��*��#}�
8Y�.�9���3Ie2����t
�H�vtj����⭴p/�z���s���iy��O%�M�:��r�} UyՆ׍L��D��K�"�L��<����,�/I�����.y:�+ly������k�JoM�v��=H�o���=�8�[�Q��U�<�n��3�(4�UO��N=�t��-PYZmDD���w^��q�I9��۩a�Y���#b�/���X�
�Y��S�K���WXto���)1�i�Q(S�:�Q���ט�@Qߡ_A��d��T�����c�6�\��f�FfJ��R��A!���tY�C�J��*��뜞��QX9��KQI���g"]ӊ���/L���+UFU���9�������پ������q��jD�5�b`Đ?=i	�շ���ю�k*3p� �lr۷-c�`�\ܟ����_N�2�LR���ը��Cp���'d�Z���pSB��(?S�pF�(Qm~_�P�����`��.���abeP;���Q��o�}�y��A�(��
}��t /VEiyo�L�� �x����G��Çe�D@Wt��'����k��I��"1WKG�����j�mC��u!���/��4p�r!�E<����J�A~�w���{U�ip��Nm��H�j�[R;r��o�!�شZ�͟vĵo��;�����!�W�:���6���������w@�(��g�I�!�]N=�\}��;��!�"|��D��lJ���?���8Fg�bÔ�z�E��r@7�r�B��m>���rQ�X�ɥ�'	���.���;
�̛C\��v�<xf�l#�D���R����[�r��g7�7g������QAh�ҡ��	mBb�lÐ&-�_�I]6��{ �/q�4�q�g�*�]e.O��������A���H6��5��i�`���J<r(0p�$�����O¹q���N%��s�Ȝ��}a8�/�B�����4��)��W8_H'k���$��<)��{�
�z�[��_�L��uq�N}�݀C 쉎{I)����WG(��>/ͅ���@���w���Om�ª�1>��p$<_�I�c@]B ص���560���������yh����ս%[:7?+O�3�)�ҭ�����o\��玝P͹,��