XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���L��\IS�	��^�p0�gu$�_�ӌ2>Hj}J�V���E��:��F8��UN�����Q��B.�p��>�����I��Z������<���!�1.���CK�`V?���)��T�8C��4-�ƚ!Vi�xY�,�L���������:�
��\� ��ɍ�Pt���i�g�e�P
u�>3?O�-F��]���~�l�y9L�� F��вk��X4�s3�n�w ��8���u�~:Te�I�-O�5��C*�p�9�N�4�����sT��l"[���0k����e`w�Ґ��cNoK �;ǆ��ui�7o��Ƅ��R��&���ڌ��c��b'�ώFr#4� �=P�L\Kk].����!v܌@DS��ϻ���l����qhp}�P�k�ڧ-�Q7ޥ�k+wnq�r(#�%R�iL�A���΢�-;�������
No�m���y�^:ԇX�
�i��>��(���2<!�v<����\��͢D��""cR@�Wg�=���ЕkIl��J��
K�]�b��߅�F��6]GieO2|�1X�x��D8��^� $KZ�i�g�-�"ˆ�8]צ����z��D(\��^{e'1�m���DM�l9��9�J��jy��XԿ:r���B��h9��Q����U��F���1�jJ~;3r	]̷��3�"�}�z�&��eGvr������C����[q���=e �@�=���:l罢�0���ΰII���e}j�,�!�`8r���XlxVHYEB    2892     bc0��)�	�;����[�A�mO:L��E�f�E�rcG�W�����s��1^��0�Q�PH��ɑfJV���'�q��MF�;�㈋@��3�g�_�_r�7x.I���W�WYu��~���b&d�ȎC��t���V���MC�d��ъe��.�����瀥SP�U􆮄p�EOPZSѲ����ʴ�ԟ��o�i�E3�)�e��ۖ���.q���;��$�~�������x���(�3�&��ܔ=����))����?�e`Rq*������~�q��uq�1$�����0.0�"wΨ�͂��j5��7������������mŬU];d�϶y��m^drE����x���j�N�T���2�xq�b=�z�8�y�P�CM�U���ط��S�����S ��ǒ��8F�]z��v�Y��%������I%x{�sux=3g?������!�J8q��V�^t������ȷ|�t�b�{�W��Q2�b4ϧ^�
�ʁz�`�V�+ӧ�!��O�!�u9��Y|�͹Z`r\t�R8L�U�S��WnK�OQ�;.b:X�ր�Ǒ�vZŁ�`N��L�w���v��I�II�t���������;Hl&�Z�ςD�+�q^�cU<��K����HU9�<��n ����	:���2�G$t?� �E����Z�°��M|�ve��gg7����0���vC}mR�>e��"��z�By��J.j��΋�Z�k���y�}7{��g�v:��XE�L=3݆G�AU�[�����٤rc�e��)׫���Ƚ|�ZK��%A`�d*r��s귎��1�q�Џ�6�K�+b�u�
�a��.��b�e<�{VqD�`�!{pnT��oE����-�]L�9�n�O�!F�}'�/���0��"�J.=;D��GL�����I�UI~���|��#?[L��;������n��@�����E��/�i� �Uz����?�ѿ������1u�/��"�"�)}FȎq�	>	��^o�h�D����=.����>��y@^�e����E�E�ϱs���@�!qǆ�����h�-���O�~�z��d���`�O�3
%��h������3��{��
G�1,���Hn���0gȇ(U���-��.�����a.��L�P7����m����}R�b	�T	�B�jǫ�l���U�p#�� Ú@��sr�X\���[���o�:f���y���ia�z�b�M!��w�����f=(K�cF?�`��x_�� >�������';�;�²v߯�����9V�:�Z�l�SuG����/̇8�c&5���D�5g���1���Q^��9T8��
�@@z/	�A�~�/��=���Gц�{ݤo���D��T։���S*I��=�_cq@~3Ό�u!L�1r[�R���0�� �T_1�(��mwi����:Y��I��'[(�,Ǐ��V��< �`��V���-�j�c[�{���M!����J��H���]�̉�e�q���0��\Q��1�E���L�龷���� �g���E`a����f�<D5��+�q��v�6��;BXsƾ�1��:8K.[��\9�zQ�\�go ٱ㥜#O%���� z�nh�)��w=֖��]�>O)u%1f�`���ݠ�\Ҷ�?��oT��`��ȏ�y\��p�}&T��ۗz\������b��xg�i������^��"��>�<�Ot̦n�W��5�/ˍ�O6ٽ3	�Yul�pI2����� �@��]X�p�)�F�u�#(�m��ɹ�2IP'�����5�qV�l�|[����>Fg��i�mB�<�r��Jse�Ż�y���
�gd���j3'��;<$�?9X�SxojStTG{�>5��ݭ���y�!ͻ��[��%�8��n̤��s�8��T�I�U��;�8���M� �]3v�&�#O*9.׳���3v�� qAu+.T��]��?�k7�-d�E���y��?��훂q0a�!�r�
�`{�}y|���������?� ��
�O��dC�8���ku�@�zL�q]�&�"�&�Q�,iR_W$�"k��5&������݁�}��GK�����&n�p���Ȳm�u��S���{��h��=aX����}�l6���� ���ξ������x�$�@t�8�-CGi{���2RC�1w��]�8[�k�"n�7��(����JS�יִH�"D�˯��L|��58w;<�k����{���x�R*zt�Q�X`E-���������)g:��xh�Gb�K �}����ŉ�E)U���.���Z�ѡ�l�nQ�8򰸠4%r^R��$�۴�Yb|v�
�W���
2��6��Xt0O������a.T7K���,0��%�}kK_����i�!B%������I��υo%U��ȩ�g̖?�^(z��pN�]_�_4z&s�o��卖��ZJ�������?�x�)J���w��U�Ӱ��Rd�!�F� �Z{��6���迂�,���5u 7��a1���/�eV�yD�Ĭ��x�A�hW�K9��ً�C�p�XM�" c-��
�
���l*?��o<ڵ?�`ʟ9 ��֍D�3��P��MP!��8�k�����|��ǁ;ԫ6�6>��<)&�'u�>m���Eڰf�	�fǗ+��V�����(�侷�p;�+����Gd��c��H!�T�D<M�4�����s�HM�:��a�_#%y���)�.��e����ߥϿ4�~S�����<����T&�¼g�'�~��X���ߊ_ xT������uR�Ab�����k�w����KjY� 
�M���|C�F��𼑡N�Y�g����0[L�Ro�(���a����c1��~�F�^�3g�F8I�lk#`g�Ʃ�V&�����v4��&�6������K��q岗�l_�Z}�z P�E�+y�@i��X#d�}�ՂGK�">3�EPUSZx���{�~WAEu�������9