XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��/��<����D�ݿf���1�S'~���Խ�fRQ-�:�1J��̥h��cZQMQ����Y�9���/[����2����Hfͥ
������q0��p�k���o{�< W�����l-�F��©nUF���P*F�XQ!�Iu N�f�,��b��p��I@��+�k�y�tɮ���*�y.����������_�!����[�vj��&���-�� m��&魍��<p{�#t��l���j��ׅ��p�}�L�d�m�rX���͕� ��cȾ��.P�����d@�t����\�;�j�
��|ɩ�r$�+���Oӆ��c�׎�uǇ�z����´$1�RXwrR~�0!y!���&m�;F˂y˔���4K܀�I�Ѵ�sy��+�o�Hv�j����a�1(�E�	ZqX�J����d9L��!��S>�O;��,.��դ�>����x%�Q'ua��-�f����Os�p��3@;��ӳ���r)̼ ��Yߤ��y��t��C���԰x�FҀ�����e�T����o�*ۈ��SG��j��1+���SQc�:i#�G�E0��e�ԗ�"i���;�cq)9h.�Z_�с8A���|ގ�9Kr���}z�r���SX����ϧ4�M�xmM���PК@�jhd��uPt}��-���(L��9}���X���B2�2Ԙ���N��=�?�GFNCNm�Dۦ;7����o��`��ӥS�:U�v�߲;���K3�VtX�!XF�XlxVHYEB    28ae     b60B��֒��)�X�*�/���̇7���X�-~�X΂c���Ԙ��³����\>�O���-��4]�7�c~�b�?��c�i�^�Z|��מk�L9�.��ϼ�+jGa'���ACK&Dq�@r �2���vb����j[r���v� Z1��aΤ.�G�`�

i*'���7��go�wP����E-ϳ:\1N�E����Zƪ�e���~�q�rr�Tl'��4-��"�"�$=�.iV5���3�V�ᒽ}��ښ��-�9�H��YWJ}���G��%0c���I�n���iݏ�N�V�S}b�m���]���� ����Ļ��2����ps,w�^��!�x{2��Frj�)2W
b��w�~wE�ί�Q���$��u�K�,�����Q�Q�_��".�̶�=Y�s]%�Hxr[�����"Ĵ �v
�vBh�
�*��PaEP��j4}��m)/���k�[�o6�f����ԫ�ZXM��Q��aGo^��C�J�+��m٘+��?��P*��sXH�c6�d��ߧq)��V��9��n|s�N�����5V9���ܺqij���~L��V� &$�7����M�`����������LzM�yb�>kј�e�L��)���/��,�(u����m�&�Sc�V�ߡw�I͂m�*8��h�\�(R�޻�J���^qW=���6�ߺ��E�M��� %H�Y��,rp�C�E'��D��g�Bꩪ�������4b��/ �a;��-�uԹx�fP �~C���i�3�w8Րij:6�m�7����.�	8a����͎HnO~��5�4�t�ݿ�|5�<�Qv�a�HW*$�Z������T���n�uz��HIh3h-�$��O��dL��/;�e���B*��{ژѷ@�}����mXJ�tq���;��M��fe>�((��CYa,\�B�'��8�k��H�j�֯ �;2�Y�!R��V� ߝD��$Ff>��h�յ�$p���=9G#�-coײI&o�5��U�����P1sX�0����
�5o>Z�v��ۢ��]>�t������i4����.�w�3�eue��S�oc" �̩�K���g��@�b��B₤�Q�Z�l�� ���g���S"tR��x�M����8�o�=
���i1�t�|����C���Ky��Ӡ�����c2�� �'����1����H�>��u�;����
WX2U��	a����5?���9 ���.���	�K�K�A���%��qxSk�Dxy��I��5������l�t��[{^�a4�]�L�ʎ�js�t�>^�p�Ϭ�a(0%4Bf�z	l�K���~�����y�A�[���@*�Gj4��i{gt��a̯��ݥML��*�	���y:���ʶD���L�I� �-����	2v���#�햊Xk���""m_8My�
|>F�mwxTl'&	��7�̛W<�������4���������qm��e�帛]H����Ɨ>4`}����A���2�-%/[|�p�x�O���?M
1������!��1���_��d�߱P��g,��
����뻋?H"��tv�QU;���I��=��vL�	��'��\`�G3p�&*�P�!�8�D�ә��Dr�j�|w1�%z�V����	�U�?������!�[���,��o�o�ZGA��p߇�C7�'s�53�����{�����:��=�A#?���H�0��ŋ�+֩�1h�c5��5U�U�[��
��7$��6�8�f�QŇ�������~J����W�//�oG� ��,�������A�ґN�� �+������;�P C�#�����ce��	�Pb��O1��9ƙ�("��M����^�L1�ށ}�� N�%nY���q���m�����+p	�>}c����m{-ZC4���F!���<,$��i�y�����~'�Nf�e��ܙ�~�TBB��o٪��2��d��3����	��
}XH�xje�?L�s�2+�O��̦�]9����W?���dD`�*S�T�h}@K�$dwZD���Re}�u<N��R���w���.R$ ��f7V��ߙE�������ן1?����yZ�����I2[�Ϸ��[��vމ�0��L�X�^�ٛ-o<��;;KNM����T<�E�l��+h?~�4�RA�pq�c�X�����э�Pe\5x�ϐ� %�A3��ן�o$3Z�W�UC*�3j�S^}N��x<e�M�lE�@�1�]�|�%�f<TGL�c>BY��l,�*�Kr�2։e�u�����g���WŤ��C�[�u ����[,.{�?��V^jJ�A�Pjt���kc}
���f5�3�īY�k~.{gi����O��:�4Q#T	%�Bڃ��Z��1�
�����T|sꔨEYxrT`}���Jj���qK�rΦ���%�^��a����H���'�����f(�I����1�I痵]O<Q�/��X���WΫ�(�&�Qau��_7���7���ٞy����4pù���9
����\"f��X$s?���.V3�v��*i����^�De?��}�C�V���/dK�;Kp7�|�y�'�������>1�X�F�Y��lT��7�@�(��t]qK?[0+�xͨ��\<�i�PQ9ѝE�<��P}�2G�O���#���j(uM�B\�j���Rl}[�H��' ��V���:�`9�ET$ O�ìN)	���h�>�ٰPg�
*v��mjY�����)�Mۜh�{����AK�,�xg�m)�J;E������*$U�k��:؀N:�xe��}%�L2O���>0+-th���F�eCs�T�tno�w;�sqp�c
ﳩ4��ڛ��