XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Y!�tv`��4��6��z��[7c6�6Ld��<!<��>�P�[Y= ����'Ыy;����<d]Yߘl�]������<#�K������<�y�Z��@��~����<V�a�%G�g��ѯE�ƫZ�r�L࢝�B Q�z�guD��ևd�Ky��E'K�&��v%����U/hs�e�h��_�H3�[�n�Y��vM=��<A'���t7LM\S�Ȯ�sR?�O�K�Z�׺�k5�E�О���.�ç{w���ˏ��࿤�%�=������!��l���Ɂg�|�@������e���Gx���i�L��WK�6`$Cs��i�Gf��t���g��n�*�Lo��1��|���F�B"�4g�wMlK��T�u��@|A���)�2���`cR�E���L4H|^�ɝ�W�%�ܬ�`Bt��=F�6�Iͺ���I���un�V�*E�#9?��&�euh#
{�_X��FV��V����qW-Æ�/�OѦ����:ˋ���1 �vP��W�Wc�fM}=��ղo2���=�#U+P�X���]V�M��C��!4�pS/�D��O��'����>^�l���&�mg��#y��l��vٜ��L>�]RGó7�)�%5�]����0��.�>��ޗ`�!�(��G�9�6ح�	QbL"3�"�}l~��{��D@�p����ɟ���De���!#�(lc�E�wy5Ay~�d]��c; �d�+�ܘ��` �J��B�E������O��!�Q��)8:�����[�^�XlxVHYEB    13ba     770�;���l��:��W�Bz!�Vp4��)I�����/����{ ߹H���&@������0ؽ���
iy� GR�S�ʦ����n~쎏�@�Xb36�h� ��'�uB-�mϮ=�Z�u�t؀^����~��+�6�!��'O��֦�z�B��4���5��A�r��wE�/j
�x�.:�������(�-Uu��	^М5F��h�$�U��Ӝ��M/`E�F��2�����,;�8�t�g��6&��9I��<��O۴�x5a���(�\�~�:Z�x�A*�-0�3$��n3^���IB�1|�>v�&�����*]�ɾv�sX{�L%_:��&L�l+�-54��.bPiDٙS�.� *H����)3�3��d6���f���L6�������z상��m��z�ro*Tx�� �d9M`D[�1��R���B�%zT�'��WO����-rMZ{+t��C,�6%���D4����@�ۜI$�HV�B�i.8��ȷ�2�B7>�~�MY(���?&�	����V�l�d6��w1�����W�QR��Ct6�����j{tO�"���<?.�h�M%��{ҬH\�)OK:�Qi7���&�P'�q�YG�	�[Y�,�^��G]ج�����R�؋T�mf������_��
�e��_].|3ɾ,�M|x�8v�pa%4���6��և6�
�J$S%��.=� e2u��O;�����L��uM=�@8z�I~����'@o�;���"��q���[��,ovG�0��$�ʶ*�\͘����4a�ՂE��h��;r�f��� ���1U�+�6��K#귀u����9|�7D�J��(�#�E5�X��DG�:�g�����|��i��+C���A֊4�~E_ɾuK�<���*�=�W�k�ȣw��2��m.<tݽ��A�F��m+��/)%�Me�����PL#T]K�W�w�TM�?S���7r6�NVڤ�ů��ZN����G�sl\E��P:����h���_;�����Z���|��L'����	���\=�����s�F��5V}q����8�ze���F�'у�[�$y[�:+C�2��ݞ�O��~���:�e�.�z#ׄ1�	]�Tn7��8�u��D�x�~nk��kUW毧����Eᅩ�G{CS@)P!uPpl�+��v5['sg1ϳ�����$�K�?�{��DNvN�0��3lWI��g9�7߃c���x���s�-LWY��v7%�:�Sg4:�9VHd�H?��9�,�pMW ��$�urV��%����b�ZFlu`Oyp���J�HZɨǧlk��
���@����?��K�aH�P^�B������$2w��\2�Y��5��ev�w��ü��9j_�M�����f2��	��OP�Br;�/�ML�����0DsK�:����3�V�Z���b����I�|N�������A�8�r��� *���(m~Rd9+���=%��'P�N�Ԧ����^R���M����e��8ҏ�������P�A2����1N�f[]8�����1�=�kU�)IO�	�U�C9ӫa����nr&{�c8kb�N��ؐ'��މ�M
��h;��� 9�L|�S5zs�2���>D�9���E�������7 ��b}���,����\N� ��(���&]�ƅ�b'?�v�)z�EY��(S;�wm����X	���d�4xp��-,:�C}
7.�(�"e�bN����H��bV�q�����m�\IX�.hOq����/���Mƨ�M���Ȍ���{�,�A�(�5���_#�J�;&�G�O���K�]>�a��j���3hM��FX&���ݫI��#N��(����'[��a�
���ڻ��V(�