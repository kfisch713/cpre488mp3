XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���c�u ���<7�캠��9x06��s�F��Eܐ7	i�}�喂[rK��ȳ���፜��E2dK'ͺ�2��u���6�Z�sf�Ƭ��y�Gbj��;e�7n�]�*�)QU���3 �3��-�=�>&�V��x�o���P��=�j"N�F�-�pQګ
Zu)_�ߌ��x�&� X՞b��`��j7�f6����J�|M}I]G��r�GF��a�x*��7َ��#tiIC��a�DW��(؍�(!�X��ot̥k��3���&����_��low�>]����YW�	]*]���>>��\�B��ߕ4�f���I
<�e�aw��J�H`�y������J&3�%�b�CJ޼�M���TUㆾ���q��$(�;WbA�zh6�c,�P?m�A@��/ɰ9�b%��jz8�3� w�{�l��V�%��4Z��y�����q[paVg/7kF�,v@w��)M��0♶�MАW����v:}M���5j�L���0�B,���$��"���-V�����P-
G	��gZ����%B�����6����d���Z�\_J�C�ze X�s�æ����NR�fj_��t�����WF�|�� 6s��7�k��\(�F2� FgS��iE�=Z�����Cő;�j���9k ��m�WL\Yf�_S'K�yݛ�Ы���P]
�e���"��S���'z||Mp;�?�Tvq�K��]X��a�.S7��@��:�����Q�qXlxVHYEB    925c    1a60��w��q"���������b�`4#A��?�u_Bq���$b��[�6�h]�Ha�F$
��qΔ y̵��p�l<�DlU�q���`ܒ�aLQ�Ď���lET삗��[�nk�@@&�S���%���LG�Ȱ�p�r�hB�.�__	�6�T�*��U�AI��+)��1�DG��hژ)'��� +w+r��"���$�xw#Kq'���ˁ����v=٨�*�G3���$�(>�冿��E!�BZ��]�-[!]��S
�+�^��é�	�7�ƫ��n%�P�..�{��v<V̑mӪ��f7R,�|�Hfq�<><�'���r����/�����U�SP���A�E7E�,��,�~�������-hf����R�Q��ٝڍx�I�j�M�'�)�8Y8 U��"Hۏ
\�N@�������m��Y�3s��� ��Ye����2*û�(����m�w�H1�&�".�����A���#�nNV�H�"`�����1�Es��Gi�)b��M���~e���vO�)�A�_�
t���"��c&�ҋDͪ���$����8[:�[�,����`K�C�@f}j�WDŪ�͕>-PM@aI�͟U����И�N�?ѕ�gu�ޞJp�ז鏾<��v8�Xa��s�5a��v��+�8�z^����8�/|�cjj�Cq"�֠Y��>F�%Y*>`*SG�{uU��i� �
�OY�?�j�6p�d��K�U%J�jY�U�
�x �e�jN	��7o.V5�v�Zr�\۽L=�=6s���|��w��[���!!_\��u���
D6d��ٕ) h��#{�I���-\�U���e��r�0��XW�A>'tX�&R���=�47_��;Mbz5#�Z�%w�,ą�����a4-��y��<�]&���k��h��%��(�Nq�}�o�<�,<��$ٞzI`����A�Fs�%��@�{���x��sϼ�������j��TQ�[z�������BG�Nl��ֿ�e�O�VO��Iݥ�q�-X(��>�"��ˊ�oH]���&�?{���pZ�.�Y4�t +�l�������D���u���C�Wf�-���E�K`�.����iFl�bỨ���T��)�,b+�@��D�R%P>4�{?��6�|�x	S� ����C����L�n	_����Hh:$�@;t��@�g	��l8����-�*L�2�OC�Ю�{����)��O��[��5�K���E�m2">|�Z���	F�Թ��-alw�;��ٱϸ>_Ug�yf�L46����h�X�Р��Xܪ��_��}ܳ}Zi���`������[X6�YF��y��:�������j�M����m@Z��\S'޲U���֢��p�9殆VQ����9�4���Q#)d�"���@��ү(�Z�'��o�ټ���.��+F�}����$����_2m��/�+�TCڸ�,��ts.裬�˱�N��m���J�5����`�L9D�H�L�T�3h��GDN�#��#����N8!��	T]HUa�g�89�h5��BZQg6�kvdx<�T�k���\�{ɂ�Q�f��2��A���!�`�o>�M��'�!��<�>�A����\5�9% &,`d�c���>�p<�zѾ�|9^���W[8�̥ >d�Uȗ��d�}!NV�Q'I��`&,=�����f-w���i�M=my6bft�����P�u���Mg��!�L.B�������'��.�?�L��F���A�`��˵j��ӝ��ce`���Cm�D���c�i��HE�ƥD:4
�߹���c��`�&�3��dw?qX�#��F"�oמ����Qý�%�{Z�8��ji��[l<�n,��%- 	'�����ӌח����)NfP�&��&��!j�Zl�a�L�E
���Q+8�W�lw�
���@�NEa�o*H
�ۚ6��G�U�-��lΑ�KWV�^�ڠn�Q 4y�4\K&�D�q�;�?�,�iF�ך>u�)����|X��9�P�:7�h��0:1�MZ=�߫`Y�Q����r�J��G���2TIү����e��N����?;�����x-=����&$i��c�����%�Y�1imM��m�=L��<�b���jA�4��z���� �m��"��t��}��_�	f��쁈ԮtsW�1�<!�NҮɒ +�P��-N6�z̴,�s��^ܝ�����������Ql���E}̳{�:�[�n��oso�k��ψ���{��s/!�*n楿BZ��~!���f��R��y�O_�hm��О>�7]�s8�hqנkJ�z3�?Q`��FX�'F|�W�_R�Ƽ�.�v�5�z�r�$� ��8(į����F(&Fp/n�҆Jl�;u%"�$���5إ�|���]n�̸i$X��v�;���!��U�,@T���"*����`�e���W�/��c�(� ��`J��!�������v�3�')!�E��{����A�T^h�^�5�R�/G�k�A�X�󟣰Z�\�˖ʔ,FC������=���ͳ�ׂ7H���W��-W1�j`���BS ʇ�Np�V�Or�D_�>x�c=;w{-�3��F�?BvbKf�A�]	AkݼCM˩�v�[��^�������xhIGZ�HF�BCxB�&�2�_�+��0lrsL�!f{�:uWvt���~��A5���"�+ǂr����.	/;���ڿ���V�V��ǔw��_�{Qc&��ΝT5���RV��b��k�;�k��_t_�&n4��bv8�����EҌ�Y��|D�5��≀2�AJ25�YJ�WO�娱k�XCJZ�A6�hrf�����-���D9j�(���$�Ac��k����**fY������c�'-�I(g^��g��o$�V�FU�}�x�5A����09�F�:W�[9�#	�A���i��A�sB�)J�}��;��d9����/*���b]�k��Q-$1&V�9��*/�I�5��	�N�ݙ��	~�y��N�C��7��3O��
YXܻp��B2KD9��~�6�MpMIn�������@`"N�ɮ���A��ڵ�J"���0K� ��)�}�.�g�{S'�Z��S@g��Z��~�G���-�Ü��0�GiF>(?^����G-$���Y�ڛ��)�^|�4�D�u�+�3�Ӄ�qyZG:5�<nh��/B� �Q���J��+���R;MB�	U޴
�!�l�܅��H7-����uDO).�Gⷤ��)AJ�T�"H�4q�+;{ɀ��E�?�U�`<K�n�j	r�t�QM��05)[q�/�Ǥ=����,�A���ԕ��-��� t�f����"��ػH��?p��G�UAV�h�a<3
��r٥�YC.��oj� �j���ްW�H�g���Z�e}�vZ2P���?p̞�+��n��0���3��6g�a��_�=�$��d�ƃ������5K'�n�� ���ᦜ��;14]d��8v-pE}��j��j>�Rě\]llH�q� ��^�o%��Pr�4�K�V�X�j���s��HeMT��� :��7|�y���2j��:�p^��oSU��ncBf!.�6�P��m�a5�Nz�ҩ�iH���ߩ���V�V6�C<*۞��`�9�pQ��Y� �����#YJ��;���+9�^�>)����$��`y*s��	ӆ|��4�Z[{�����=�Wb���p!���ù��R�Q�䝼&H��
������]{��G9�`�op�Gr�B������<��r���Ն�f:���6���˧#��t0��[k�e��~��-���(��:���zp匫I���4��.�l�)�L&!��ڸ�ѺBe����)��������L8��w�~�z�N3�+V�O*�}���䟘g
ek]��N H�*%�7�"(�ؼ�u��;�3T��[�*�Z�mA�'[t�	ʊu�ؚZ��0#r�l�)�"��rR3����]I�5�6��ht�쑢pN�ɍo�jk-��x5����7�ᥥ��̷hb����E�^B�M.����'��[�3כ�-|�X���1,�J�r��k����\�F��S�*���fy�ł�����_ ��	�5W#i����w%{=V^>:K�9�N|
���$v��ĭ>M�K��+H�ow��_'�2[:K�tx��9���SԼ9/b����E�-�r���d��m.x��v�}��Z��җ�߫�<���>9S1 ��~U��|T`�w6�e�8aTW����X\-�i/�v�ˬ;*�vC�vEd�;o��͔K�@j$m1R=�����̺�A*�֋��P�I�T�����5]W�	�K������H�^�(�Z�T,%]h*
;�g��u��7����fEt�]�q�"�~�Z�G��������*����N�X8��ᅥ���~�H5���:x�
!�b�H����5b�߃�oh��1��6{	��<�iP��K�X��ŋ�9I������}Mƺ�a���I�Ρe�$���s�+8��ٶߩ�eaU��<,|�Yd�Jm������#8���L8$_.imƬ��Ml��g޴a�e� ��N��w�(J�� 
��;�^��4*s��M���b�z'�Z���mFذ�j��]w�����S޴9��t0V�q�h3�p�̌�уQ>��{�%cv�+��G�̇�x�9c2�}���%��"��'�� ��+v�[���͎�F�:t#����uP��{c!�;߂�w�|Wj�3�P hZhu�3}L�AE+I���_N;}�~m���uu������0s�~dl�u9Z�Ybm�d�&xH0�d0�㶫���C>}��ҳ�c����Z��h����N���I,�]�B"���GϢ���y�B��G�g�<H����	�`�B8�^���p
2C\ti���2f��,�-ğ!�l?H�e9,f.��ͻ���l���+ef'����3��RJ�q��w}��,-\�v.����˺v�VT|���rjh�oK��\/��	mԝ�$�&mt+�R��<jj@nhj!�7P���b�d�]���C�7�ԩ�NѿĐCcb���x�����(�}��O�����X��q�0놚��37�?|�!Ƌd�`)�!<}*�f�gԹ�ʪ�zxpv��4#����?L��O�|�������>�FYC/'�v�ͷ�+Mi�����t�aU����#"�L�_���
�VZP���)�ة���J߅Q�nQc֍s\��<�!�;�U.�1��#�sH Qh[ ɢ�S�F�� �;��6����
T���Wm�����}��4P�j��K6�>�$\����x�+A�Rw}V`Uq7���!>��o�o����q�����Sȯ�g';I����Qu���[Ma2
���L?0�����oSqՕ�޽�w�Q���"BJ�𫱋�m���mlO�j�=^��E6&"n�����OL��b����nl�縖�噫�b.:���42��{�`FQ�9vN0��>�8Yng"�VF@��s����ҟ7kN8o�g>1��.N>p]���\'�3����t�`����؋	��j�c9d� D;��l�_�m�-;wH��։&�~�.R[�?��E8����`NMX�u�78��El����W�7HT�8��p3��I� n�-���?�>�ѓ�>��ؔ��:^dV�.H�f�+U��J�5���<=	 ���0�+i�W�8�D'����%:�2�ܕs��	���c����:��!8�q.=��~�a�k��'%Αz��pLd@��Ң�U�!�Y��2Bh�``E��iL:���S�{㋐�ب���3S����o�%8����OPe�s*�-�A�]��E��^�����c:5�
�ܾgEDL�������dxq-$Pa�$��Q�v���\}�,;F�����F�漾r�A����2=�tlk��c>��vv���|���9��ATSz���BV�P�~%>���~�L����e����[���Ȥ�ѝP+.�?*W��VÄ�c�+.U�̴��V�[f'���u�m㨆/��|/��6��ύ� >Q�4~��vO�5QC~31C7�����N|J��z�gE�F1>s�%�'�X����/�z��U�u�^�"tO�9̅�V�YK%P���0���H7�X�#��Č$ �����[�D�vR;1�X�8a��_��z��7%��n�(3H%J6Ms��|�K��Px�,5��&��y+<�	w�e�xB@�≝�&��N9{"��ָ�~e}��T�>������0B3��b�M.=��?��\�\k�7 N~���}ꖟ���\ܚ���I��۠X��p$e�NGȟ#���L�֍s��zD�rQ��$���vg�����F�� ��S.{�4ϸ�������FOW%�#</AEG��< ��}̄1b��^E*t�o���q��Ģ�Y��Lp�K��.EY�+��)2g��X\*�;�Rǫ��R�ŉɸм�*[ �u�[I'{k�#�4���\\Z-q_���0k�%���۵��7�H��������^�?��qP�4]�Q�}��׶���Hy��~��9��������M�������k7�( ��҂1[)i1E�n^'�P=��$�ٯ���$�������pƬo�͙x? B