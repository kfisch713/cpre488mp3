XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��������x��M���AJߗ��!�+�N4�p�3ZK�J����;J|,U��A�b�4�(�.�b�켹4�窊��0�(�j��82D0sN�z�X���L�`�7�?]z����,WU�-� �T;V��~;%qdR�h��n�L�r��Bڏ��8G�K-�!<�x A�Y�s��_��z��&ߌ��m���`m3��	i��\���өbvF;�j���v?��qT���w>���i��J"b"F�(�f^c�G��<��pY��U�؜ޔ?N��>]R{M#��rR�P�\�N�ȩGر�U1���2�:/���F�{�D�Av�5jzeB�3��z�Xo�@�'�e	�q�/�� �N	�� Q���t����"�)G��_��'����ܢQeT��٤[U���^[�4TA�X��*�28y��AJ�x�;�C�ke~F�J&��f՚��\2�>.J@��3��
��(�{��'S3̎Pw�S��K�_t����>���n<~I����U</�aXk�h���(�s�j�����J�b����	R�rқ������.2#Lz��'�v��N���Q�Gc��C��l�R�T9T��e,1��s�B]ݨ�al��*���8WRM����i�x=6���)�A
7m\ꦑ�06�A!<�F���M�g�ckة��(v�J�q��6����rޙ��=+�7E1P��7Ԭ�S�m�d��jN�@R�c�MO���F��
-Zq"�3�D�Nh���8l��7XlxVHYEB     f9d     6c0f��ⱦ�t�YL������ x;�ѯ�0hN{<��q���P�~W���]�
�X<�Fb�%���9�5�"M�}E�8�ќ#��^���B{wu�7�?!lz��3�B�9D����;�G1W�\����8�RҀ��Fz��s��k�I˙�%�E�p��k���EF�̀H����6u����7Z�F�;��>~EO��:/��OgX� A$�kL|�Ŕ����` ��3�:�s�+�H�ǌ��� �u�	���u`�B�s��
~;'�n$b�;J���=�vN���pf$5wPb��Z(f ��7e��&A���[s Z�
O?�3�7r3�Ű-f���xtF� s�G���1������i.ۑK�$��3��o�S�����+/V	���|0�� \FĿ��TK1B݉�(�١��㣭}��`s�%~��-%�ӠԘ5"{��u^F*Sf �X�f�����q��D��U%����y����	=����T�ɴ���E�
%Yi�(g�[2G�c���+I:Ǜ즼n�3C@�l�(���^f}Cym�ͅh��?n)+�[H�!~5?��YW�~'k�u~;L�2��Ȓ��Ʋ����ar	 |�;��I���Z�-�}��.�� &n��ΣF���Cv�����P�\��02v�D�e]"��j�iK[#ֱ@i DS� 4��B,�s3,j��M.�8�����L����wmNW���Bǲ�ԛ~9�3�]:0��r̷�f/ o���]I�ig	���D�}��p��Z�p�E��w1�̑i�k-K�P���������C헃oݵ1�]�?���������'ٸt�1G��a����Qa�̎GIVA7�V�߄�6�+"ZT�>p"�z1�~%
�c�;D����5u����d���#�3ɸ��~�F��� �X��o�6�to9)x fM*�'ǭ��A1]�g�M h�ZY�6^��žu�((�����)��(j9b'T�M%7�T~ RR�
 b�0��]u�� ӌ�!@a�:��J�}�����a�T�l�ˋ9�C�L>CΏ������M�D<��Z(�=9��H��B�s�TҸۺ0�'L��o+�d)ݽQ�3bszg��p�,�x��h����>>E-x�;EK7�,��8�RP.]O���R��K�Ά�-�)	��ہd��^'q�bZ_b�`I�~�h�������	���j:ɓ��BM������C.��=���l�[����i�+����]5�F�'Q!���jk�ї�xh�ҽ䵆� �[��i�����Z�?(��eWR���.�Vi7�cX����t��Y����#���BL`}	]W�Lƭ蚻�¬�>��q������j�}��N8��\I�k�@�U=I�?�P�xU����`9#��7P��:6k�[t29��58��OUIc��7>��b��i��rC	fE���t'����&ڎQfyj���ԧ L���Z1#��I,�Y)Bm�U�A���4��~����l�rAɳE�Z~�K=Xˁ��_�u
�h�zÐ�8�$��&BE�d��Y�I,�
��
�d���4.�1�jj�!J�"����ԉ��>g9
�drWM��Lj=�G��1`���X�$��j�G�T�eD�b��K�
6!�9L�g�3I���#7���s��\X}\ �C�
�r��X���Q}��cG��_��g+�hX|�<d�Q#�7�wT�Iȏs+��6i