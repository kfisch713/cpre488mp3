XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd���[�u�!��ޙ��zÖ�������\屒�H�L,4�����uߟ��#ē0�{5��ei>c&�PhcA�{hy��"�\J_͑b��or�n���A�``�ǈ�-�ۡE��l��QIθc�ZJW9�8c+�}��$��2t��Qё˕3A�"v�u�ɆC�h���K}X`߽1�v�8��٤.�ȯK~��JN|lD���R�)�C�n|�M�n��tN��%�U-�M���}n�?8��\����n�^L
Gs�����ê�O�|�Л��Sɯ?r+��b�E�@M��M/G��rr-?&׿
�VTA�6�h�)�Nyj��R��Gw�s��A5�÷�1�+Zb�X���m9lF��#尮v	I\A�CB� �*��q����l����Ad��;u2�[n��wbX%2��ӯ�����lV��f�Ze}��vi��gB��? !Ϥ��S=j��Y^Yo�ԉ�ˑ��A�T1EekCq�:=5& �h d�>��M[�i��k� ��1fM����Oh��\�mm�jG���WO���2�V:w�U���3�۩mA��5/��Ï��,	�b��[�r���Y����#�������=�Go{-p�d~�&OLNn�H
Fu�
*�ݦe3G�GH�5m%3B�~QB@ŀg�ͳvM��s�B�5���d��/��􋲊f!_��n�Nle�+`�á���ŕh@!�7�@��9��,p�F<?g�G��ׯ�<�M�#�>؎?�V�.E�Tw�˰XlxVHYEB    5d54    14e0I�#h���U���B;r��5�
��H�8��r;���}��'�a{�g�ʶ_������ޝ�q-+����/C����g�1�Y�
��R3C�wMeB=��K�,�ކ��|r�GHG���>�@[ j�<��+8�,�ꦸW�P�HbGw˻Ż��b�S	B�rЍ�����86Fb�� _VZ�dfu��jF�(G%dy�W߽X� ����g�w���=2�<>gڢހ��=����Q�üe��aGڌԃ	�F�]���=��zƠ#8��)ț��A���:XC�M��t�,N�ٶOL���<�ǝO���9iUm�hP̹��v�����hl�N:��үi�cD1�����.��αr��ﱴ6�g�4�HS����R��VM)��J��o>89���8�K�����rvϴ�d�t���)� ����e\<S������ �s���2�D*�ӽ���s�d��uu���~�ؽf����S�bҲ����pa^�A��	[ϴB�`�Kn���X�/�D�y���=q&3���ORw�Nޜ��(D@�n�2�r��ua��ǌ4��7�ފ&?�@d��9Y�1_A.)�E�k%~����?R�Y��L�ū�
JWHМ�v�9����z������f�s}'���ޤ������Id������)�d��=q�T���;̷�<�"֧��C�'÷�+��+Q�_��S$�Q"�R�����Ѡּ���.�l�h�xk��8	��k�"��f�y ���pg�쭚xj[X�L5lȪ-�NJ�<�#��Gi��n� �(7X��:Eh�/9���	;C!�%�Ԭsr(J���'1(SQb:c-�Y>�R^EXD������Y@��=���@)]㌄X�����^��$���cY4�dQ��/�΄P�� �E:e��ۨ�~v�QlW��yp�tZ?c������"��2S��׫��J#�ʵ잻�?���Y�.'W�� }n4`�ǭe����	W.é�R��	��P���s�"���\"��Ы��L?7O��cG9o���Ȕ5t�Ӫӡ5"	��e�B3��b�MU�?�PM��؊��S��|�<I<�}����a��!-tR�-CF��;�e*�i(]�6�d��7��[b]@�͹T�u`��Ϥ�b�)�p|&c�L#��g4�����(�'h��V�^���Ó������Cp7�\ ��5ܛ)^~n�!��L~Ǿ\6
d/��^+���Xz((�ߒ80�;.�S���bCZ����F��' R��,C ��1C��A�SW�G��(���,����h&R���2�_f��4�b=II,E�	�2.;"�� Ē�*
Q!6���Y��Y���f	��xk�.�ӐMo8� )��ۣ�Dĵc��/��A:K�uө�*OJI�5V�Й��ە�B�q O=�@�[�Z�X�9 嗪}a�W�g�� 7�J�P��j��&م@{Am�P'Fg�Q�a�D#������eB��jK F��ERp������iP(Ds'
7��aJ��X�x�#��n��9���$'@j!��"�Ƞ���_�KVl��!o& 4|`��":�O}U�ڞ�r��F�ew���
ȿ�Y�Jԅ��Ⴝh��*�W��l/$$��`�J¦uR$�e��h��0������ĉ�t�3�-azh�7#�Ӄ�S���6�k��j>`��5�<�+��q�>�O�&&��o�B|\7����Fr��{y�M��������w�]ڦN�=�%9�2�p�,�Ju2wZ�m˶�2����tW셗��o���q�t��r7/)5����1S����߾ ��Թv�>f���"��lz�/;P��&q��}y!^z��*ϓ{�t��M�6�������e���߷8��L,ԐYT�\�#�8�L�4ј"��(�zO�$�6��@s
�+��ŠNL ��W��d|u�k��u�o���ʏڌ�`������%��~j��ҋ�pͷ��ۧ�����y�mLX�@h�G݃Y��1e����C�b���kޕ�?�n���|��ڻ7)�F�}Y����c���)���>n�E	�A6Y#��ś@�1�!JD���q�
���	ذE�33tu�=vN��/���._��m��<!��v!�,�#%���=$~U��yiԑ@��hZi7ba�DU�����{)TL� 0Nzl��2X�yRĮX�F]~�6<ߋ\�o6���Z$y� T��m��)�0�+��Y�}"���?]t<���T:S�:�W��]��b�bK !�sucB������X� ;��U��Ѐ�Y��� 7�܊���k}Xݐ���QҮ�U���pF퉿*2�)����,uGv4f���r�ɍ��!�����"��B�Oc~�bw'>j�����ggĮ@���*�O�����J[m{����2{���>7���7M��+�n�,�%�7_����?�EW�'`���'$���+:��
�A|���
�0��%������D�0�ߓ��N펡���ΦW��y��� }����df3�H�:�JW_��|ޕ���9ci�-~=Vt�h�����@B`mS�}�vj�S�� ��;Wp���x��N	��{_�q�l��˵q0_ƿ_�[-b�x~��:&�Qq�	i�M�S��8���*j<dɵx8��J����$�	�-�v���~2Ϳ��¨�HT�L��+�lؓ�+�(#a�)�3c�Ts'�u��#���_�P�p������XN0ȳ[�qjp�r��*�`�v�%�&���ޑ�3�}jHx�I��R�xn�\�jXim�.>�f&u���5�f�-�m����X�X������X�,�ׅ�I�<��{N ���F�F��,�o\\���B��V'PB�u�������*��.g�H���X˜�����ݝD�0�����<� �m7Ѫ�X�N��M�m�����J�W0�pn��ت[��vw�F��-����R����[6��@M��F#��R#���z*I��^���q=B�7�M]#�������~j׺��x��L�.�s�ŉ�1��^�J�+�R�u����m��@��)��4�$<iP��t�P������x-��#��i�-�����/r�
J����S[�
�
�BwN�����	+�ɥq5�X�vw9Vb"���=Hh����+~B��ݒ��Z��9��x��sSX��ğ&\���)��@����h��T�|�$$U�R$U7���v#��s�G��w�Ӟ��%�2N���i��	�N^	o��J��'Ϝϗ����$��h⭇�k��`��#�!^'��G��_f���ӹ�k�G$�.���j�����Qc�	�(�
��U� ��l�S��]6-u����9�ǒ�2���^a|�в3�w��чz"��Q۽������9�A�zx�u�܉��
�l"q��I�[�����K��3�y���c����&M�#����(�����Ñ.�
���=��s1�+�U�%��pZ��2VP=�9As(2��lq����.zx����\g��H-��%�ńr��v�Ō�|Zj4#�\�Y﨤�<�UF4�2��h�$oG=l���H�$�W�.y���ga����
*���+L���U�z��r|���x}#E�������oe�Ǻ�V���y<j%�'Uv +��<'�b�{���� ��%~=��Ζ�i~�N�ID��B�`��R{?�m���as|��`e���+ɔ-(�jC	M0�k|�d�*�,e7' ~{uj���W��>'v�x��~�f}[}|�j�ң�l��V��*&�������cC��q��5B)�'���xde��Ҁ��R�ʨ���Ӊ\jq�p�P�&?��h�W�Q=�P��T��P��|>]�ۜ��}��JOoח�,��%��F�o��?�����{�g=w,�4k�4�Ζ�3U�1��ZM����vI���֛s���ϟ�i��g^�淼�C�O�iq��L�H��u�K忄��:�i3��y���u���(�`��l��1{kWɘ�U^	�m��.�K�
T~sR6
	�rW���-?���Ɵ|E��G��\�W�g_
M���Å�H�	R�\��������8Q�qY�mn����8c�+��_�M��+|	R�����E�Gzz!~2�����P�$V.���P�(�L>��Y�#a�jT7�Ov�}����=�/��0���C�4 ho=�g{)gk8��1Ν�ނ�"��V���?h�\Y_p���)��?K� �2�4����I������Π�&���m���m�/�&�(5��4���b��Z]Z�cT�m�m�xoV���=�qnQ�
��ϑ1�J�,?���B��a��Jc�g�r�,��꿯"9^SA��.H���yj�p�`4�
fO�w��Ɗ\��ޫ�:^�ʠ�jύ�Y��y�!��sතs���Q�"h�Gn�SL�1�ey����\j+_�r��G�>1c�s/4�����0(#�߾�^��Se4Ь'K���_�w��b��Ư��F��[�*kYȌ�|Fx�!"*T۩�`B�V�2�%?{߹���
r^�1���Z��K��e����	���{��G�8/.$�fcV��#PUP�����M�����L���S����Z�@E^����L1xB��< 2Y�<�b�d'��\z�lyD� |^�L�o�����9�_|?�eG�.|�E�!^�h�n�#�Cr�nH���O_���������\�V�yu�#0!cȕ���e�����5�6���+�xt��+�/��^k耸��|�pc��$��p�D��u�dh
�&�u���l=��QW��o�1"�Y�
R��0o�6���~oͷo:��p
����@_q�9�Nw�ыi6D���LU�) ��J^��Ie�M`~r��P�����C��@?Q���^�0��r�!h�*��Y��S�9Cs�a&[�Y�Jf�dC��^�
c�%�����w�m�m���"hE5lx�P$i
$*~�lF�,�V�-#��p��|�L�am���V���S�.43�x��Ӹ�,���P��	j�O;���a�l�6���m��sUږ{�!kgST5�� ��ix.#��ԓ��D/Lo�@��vJ?�I*�#��q�?�Ag�S�K����'�jM�5H�ZCW6��#�PQUh��Čb�l�ށ��K.�������������s��۠�߈��s#������W���+u?.r�}�'��R6W��h�#k�f�
ՙ!��k��A���i�WS