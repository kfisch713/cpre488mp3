XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��WOR����)�d��a���: ���\>BB�3�r(�s>C�-���L�Kf+x�0V�F	
�Lƛ�~=�x��J{�3Qe�t�O�n�i�6��[SF���} �'~4h��*+�Xi_��R]�%B?[�}�j:#�﹒3B��˙L@cu M ��IYq�u]<U��������]j�Š�(?�:��:��
���1� lZ^G����X�U8���5~<�-���H�)x|��ˉ�+&K?w��+��:u���2s0yx�>�y�=���c����<ݖ��"Y-�+C��#4K�uǴyT�u�\C��U%w|\�E�:U��1����|'շ��:`z�)�U�}�Y���Dg"p-�?����++nS���m����.��q�,�e��1�n\�3����-ıd����N��5WQY����;�rgp�B��t��Q��҄
Ve
ḅ!���עk��!��-°	_�
�0k8чAꖿ�sF�4��T�#94|w�x*�-
�߃���Ъ&�]5���p��U�r�	y�;�ْ�G�(�C�3ۇ��.��E��[CL.O:V��ӑu�<����3@��0fmU�2t���eψ���W���ŐZ^Y�[B��VE�e���TԌ��M}�
�V��X��~c��}���	?�������	���-vo�D�˧c`ȲDT�n��L�rz/�2��44�ɱC ~2lк�팆xG��qwe���	���*Di#k�ō_��g�%%��J��[�~�g�n���a`�˔G�k��e��ɂ�	��XlxVHYEB    2b75     cd0�O��b�X�x��SP�&����x4K�,w`t�8�6��l$����g)��2��T��.v1*(�71 ow���'sЦ��L���hL7;�2t�,7/a�XBY��5�{��q�9:�Q�q�[p���d쁥}�im˒�0��K��7��Lg{Ĝ�6����yX��y��4�E���l�3��?�����[���0m,c� �ƕ�IZ�@v�oJE�
(es�e�y]v�)8>�jŵ���� ��G9]Q~,c�0�)ծ������R�dKK�&B���9�Χάk��/��7�a��eA�|3�La�w�!
.*�E�)��fF���Rdl6±��9>B��=ќ�3xx�wT[�,�-��F2
G��T�8s���"�L����&��4O֒&2l>ׯ���n\Wnw �����B��
�&�;8��+b�&g�0{1+�^m_]x�i���%Y\q��3��(]�����o��?�U���Di������v�*ɍ.o��69�|���U���Ύu���F�&���7p�n�|�����%s�$�2G����j]NLc���Ā*t��Hw������LRȇ��E�i[i^�X���Ձ�ぜ�������[��m��1�.B
FI��_�CjǄ`�O67���dR�UA2Aô8ɏ��%Ӏ4&���mw��Z�پ(>[�œN��W*x�1�hc�~��[D�W򘏠fS����s�DuM���G�'.Rώ�|�߃�"������fv���[�� G�sׇ`���W�6(���x�zL��0*�˵�L/i����������8f�A�,d�V_:Z#��{*�$4�����ZcbF�R�
�ȇ����і�I��P�5Q&c�(�����5�d����iRH��r�K~�hX��Z�˿G�<@d}+7�B��ޕ��4�����*�R�0j�`�8��D�4$Q +q����%X�8�Q����A��%J�$�q<�J�c���[{'��1B��2��|U&$�7�� _eoMdZ����ι/���8��u���q�1i��$ɛ�P�]k�}������k�	Vsآ�~���u��ᶊE���� �?��p~��jVOb��]�م
�5{<�\��:�g8O�3��_�J���ֻ��)u|�@0���,����L���+yia#�8��owkꖸ#�)�\3��9O��� װ'<&���6J���-�(���,��B�	W~��cY�<��G��F5�_ݙ����������W���/b�R��G$ԟ��[�=7K2��O�z2�]���ﬗ)1w@�;Qy�p���:W��z��kQ�`���f���O,�8�e|\��~����5�($[
8�I�?(�֥p��̉����շ1���hEhk9�Ѵ���,?�<���(�:�2��fb&�E�� �9wъA�>�AoF�P��L7XZ5��B�ƒBwS�ޑ�ء�����/g��g�PvP;B�b,<���P���T��K�8��_��:��9��x�����@��f���B��)��Vah� _�eg�piz� i���k��Q�!sh4��&ɂ��>U�,c�4��BE��l��G�3�Gy~���`��mu�g�b�LT�,���C�TB Y��Z����Y�51k������n,�pb��s�&��_���[�Mt��X�0�5�4s^�Dr
:�Kx�����C�t��=�=��^��GK���m�qXa�w����\pY�v��4	>��Ʌ�#���he
%ZK���^��lT�`�/��P���҃�+�?_�:���(��?X��E��7���W�� Ub3@���F?�9�>��Ra�~1�JsB/��-Le���p䩶�ra#il�C6�\�vr4�SG�+�,���ۮ���BK���<�{��s�6���w�q4F��}װ���Pi�����I����n1�zk��� #$�/���/_q��4�s��y���T-{j3\��z�F�K��:�:��0�1�m�BN��E�|A�1�+zΆ�¯ɣ�o��� 5�|d�m�@����d}���J")����($���ū�GM�Z�ꝯ7F2��8ol��B����S'����V���(���`�d��6g���S��ro#�ɦ�ν�Z�2��U>������� �+�*����]5?q�%�AB4�l��$��jH48Ц����Qp����a֎��w��_�џ����{>0�2�G�ﰍ�K\Z�V���S\3���"�8�[��j�H�_cX����)���=g��-�1"�iaR֭;�v��xl����f��K��
H����?�l�� �.���Y��ӷ�"7���W�P��r�kj̫���ưϪ�*�q>�U<f�=-�e���G�n�%��D�N6�K5DZ�A�ޙ��a1F�4����Z,�9M:��ԫ�tt�.u�QѠ&y佒��u�ԅ��M�;f9���f�N�d���b,l����f���E�8rp� S��� �U\������-X�Ժt�$���T��_ͱ20JŹ�f�:EC2�>E޲[����Du�)���U~��1_p<�~ae�A�8х�ɠu4%���V%�q!+�
yK�C�4���`��\��x$�pQ.���V�i��Ql��	������ᶟ"�
 �@e�K��༛���������X������=R�<7�W�v�5�LO���:�^4�d�=@���Iδ�Hq�:Ү@*�]�l�t�k)e����e�Vr�(�Q1��ޅ���������k$g�H�M���b��<����ms�Ó����%;K�ﱠ�b�
�)ZV�����8S��p��l+]%���l�tYd�b���ȍ�&�o�i�
�.0y�+Z[�;{�����TV�_�t��:Z�k9`�boCO�J��;�?4#Ƥ�٩�茣0��qa�>���R�7�1U<\�_�7��Gihd�w��&�B�����^�;��:|T������7���f��4�^�]cQF>L�ϓ6��y�Cv�T{X�����%ź��s��i�3o��Y4��14zp,btA_�,gv����ˍ� s�4��DBD}�i�@i%�@i����}���jN�84A���;�@Ʒc@�:�:2�)�J��������z�Ӊ��_�S�������弚^�H�-��A-���A
̻��D�z2V�1W1�� �篫
IQ��嗊��gP�V���Q4;�p��,?��2I9��ਿ1��