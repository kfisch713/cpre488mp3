XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd�����i}s
�(r����LoM�È�J!��M]G_5/�!"R|ES����J�z��sK&D]��F� F�5�s�y�}�)�n��`g�K�5��f�s��K�i�Kh8��	�K�w�G�P1H�ϖ^�.�O?�)�?�8�u�3��ه�Z.��&F���>����:kx�X�=ѯ��f�Q���@�/��.YdӽdG�4m���	Zf\����?G1"R3�0N�.�4����&���A��n}ǲ��YfD�$ZTR��}vh�ֶ�ڂ�[0�l��y��4ަ�}��7W�7��G��2��C#g����n!��
�_�Wl[���@e\���vw���!�V�|x��̡�����vgjM�]#0�����A}4q�V^�g.�m_�1���.+8R�E���A߰�������3�y��Q�է�1���0a����z���Y�ZwD�瓚j��֏n0'�ZU/P��(w�[��$�%��+�sB�{d�N�:�i��J��T:$�>ieG3L<��_O�G�.8.��n�A���f9T��T�UIى(\����e��)@F8ι)o�IH��uq���]Rl�P��UA͘Vb���7�N�.TA�� e��K��v�xWDO�iF8b��RwGkv��f��K�γI��S0'�������rg���]}h��b���uzf��g�z�
��Y� g��&�:�9�͸�и��������
\��`2���M��(o-UC����XlxVHYEB    1a2e     8b0]�%Pp(�η0<����ܛz]�K�����je��&��8|}7����ɀ�%���O�Y/�n�Y�H4Vw��#e��kj/�O�������e}�S�
g��U���1>�q���sԦ^Qh����}��m��ZL�F<d��/B����ͧ?�����o�>������@en�B��;�M�U����8�j7�#��jw�R����OD��UK8����v��h�!��h	bӒ�fp�}�>��g�qMX?F�K2�{����*�Ϊ�f�0�wy{�'�1����Z�@��+vw�*���%l��u?�ݚ#M�\:ȁ���e⁄�\Hްe$%�ڴ�7]F���!�}*E�-p�g�#\�h��q�K�k�������c�?縓 �z!�v$�:Lm�7 i��dwRi�p�#$���W,Or��lCQ?Q�q���0ʸ̴<�Z	�3�༭��'𕮧��82��T��҂�������eL�c��;0N?w<,Ih��V2G�i�[nd�)��/� �����N���(��9�U��&��ό��a���RЉWEFr�*�_���g�
����5���+D�Xt�t���[*0��H��R��x/�E�F�.t!q���<�BJ@��l.�����ѷKk�x(�ƴo���ƍe>��U��,Y�~����R��L����o�=�?�9XSg��].��Z�s^3xTZ����!��׾b�Z��Z�i��i��������g vJ��G^�?U_Xp�B�o���/dpt~[���v�J؝�����r��K�$$�\�u�j�Y:V���q���N���J��.���n���#/.�v��Oü��{3C�4��$�Xv����}�$�9Z}�O�-�eԣt{!���GV�.l���Ϡ�ל��������HY��}qrp�L��V`�j�C +e��(�(�\9}ʓ��q����t�.� X�W��@��6^*~���W�s���1�L;O>!~���t��W�K@�������U~�4�o�H��Ga�	f!�����,����ԫ}�P����4Ş����lc��q?;�� j�(4!�F�F9HT��*����D�K�_�1w��ɻ�g��M*<��Ӫ�k�NÎv�]Z�� ���cK���X$&����u���5��M�����΢�ar���Un��RξP�ac9%�J:�հ�u�+i�{��`���6rٝK�p�xGۜ��~� �PX�8��_%�9܅�(���D���hMˇ���x�Q�J-�������Г~���1��d+�"�گ�n%:F�_@7��?�:K=�e���j�w=�v�|<�T���h`�.	�?,��#SSV�t!��M�FM;|,�鐌H��9ߋ%�@�2�G����'ڥ�4<p�;�i��`��?�2"�$���e�Oq�+�:��V:0��9�l'��j�A�~a|4�!7'����R�@Bg���ٞ���Pa&oq:��s��=�����l���Y��*�z봭���~a�G`��*���C�!��6�^�v�n�l�����Z����>����l++�E\�z���;j�0�M^ط2y	:d��5��.��*�2�;5?{��D�G���=<��DQ�R �j�X��ֳe0l2�W���1�)�LwF���>;�
�
r���޺5�c��ю�f=^B��=^�)��,�U�ص`~�Њ��7�g=��j3�iT	p�T����<�b��պ�i6�r)g�_)E���<@���nXiq8�y��	m�n
?X�od�T������B���A	R�v�|/r����^{����e�{q��J�7���m�w���$��JM��>�h���E����J��8w��蕗n�sB�'�����U����@~����e� ��N��=X��+����sp�4�Bh�6��!�u�vN[���;�A���M���+�+�H�p�P�=.	T:.\%?��h_�~�4O����B#!�v��{v��U��6v�<�5v���C�(|�֋z���B�L���E�rA݊(͵Ѹ2zUN'警Y�:׌S����QIA��,�!ux =v_Ԝ[���1����R-ו�D��U�jT�S��#o�Vc�u�R
[���0��.�~�#����D�f��*�;SO�Wr�y��L8@Z��#N1U�U�H�'�Wlk���&�1�b�}�Gm Y�gd�%�-٫�̓	-�)c*����