XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��p��Lg�/��i�d/� �`$#O��:�n@������+C��p�j�M�ƪ>�0����"q�ܬ���q9�Z�W��J���?S`��=�o��E���UF�B�^匼�:b>ʍ�����W$��5��Y<��Q[ 2&�)M�Fe�Y~��X
S�@��C�l�FO�s�_���k�G�|��י9�`5z��2`;��#0�J)��b8�=�����ʣ$��Ϧ*�����i��US��*a��=�8�e���%��~��r}9Q���y{�l ��Px��Ƞ~���a��h�e��������\�u��Qe��9�Kg�l��6I���(������2��׶2֔���G��x�fn��R\,v6J��	�[�k�	���\�8�J-{f�B��뺉��^
�70v�n��W�f*���f,�Q.��*����em�,��&x���R�~���H��F���0w��n�G�l�YF� BZ�%�C�]�����q:�b!˹J��V�m�`2��
���^#n�s��g��#-{HO��~�����)ׄ�Sq�/ZcSG�/�����ɪd�I���~�[,3Jy�t)=
��]s�1	֔ğ}~�\38_���z��c��^-)��>������Dr�.O�a�I�8�w�3�T	�����h��W-Ԑ
��P���U˕��y9_L0���c(,��jEX��3gHG^��(/ Ӥ�.R	+�zv{Ǜ�>*���ɿO� 4�yK�Ò�| �XlxVHYEB    15b2     890�o�!�&4)��-ETD�\�u���z�8U�M�b$t��Jٲ��KH�{�Ha\-��w���oB�,Q
i���H�^(�	�%��w�z4|���Y���Qk؊��l@�M��|�8MM��`�"_����0�PI8��g��؊%�G�8��DPj۞�8H�_� p��8H��Z�m���n����Ba���Q��Q��גl�=JA�y�3�l3U�E"�i���ކoy(��M�0OK�U��tt��j%Oc��>�����\�8��W��ͬ����H�rbG۰�@��&�+Q}��!�v�@a��`ǆ��-sa4��I�}�6#>gu�66���Uą�t��)���fLOvMD=��J�nhR��~��
n�����v�,*�� a0���?�Sp��K'D5�%�f�F����(�#!���*v'r�(�䵧P�b��^�ߓ��)��Sl�&uFK�ұ�;?����f`���A�� p@��0��*>K�� �*�1h�d�	Z��g2%�f��BN��ac �vO��浈�,[a�=�
�ѧ��: ���}�9c Uw��"��۲��wQ���c�9y�8�A�%	��1�~ �@r��C[�ͤ��6��R{��
R��Ր�h,�g౯P�}�М�w���f�j�����j#y��f�Py'�qW�7�K�(�j�A�v�r����;��]��W_�7*�(G5VZIi���E!w�6��L3���`�"ٜ�9h���{���-������Fz�'C���	�y�m�Z8dF����[0n�)��j;�
��Z~*�/j����:\�[�X{>�4Q��f�)1�*��u(R(��'�p�j��fMq��[�����)I��|�T��xӋ�5���R[�X���L@+�A:�L_E�2&�ߢ�b��*���.&��~�+�=�)	=��z<�Јn}��y3�5%g�����Z8ނ�o���2�ס�"��;Dh��P�Vo�W����ϥ�7X3�t(ƧG3���=7��,��D���Ķ�l�{\� ހ�O9�G�?iYsԪ������#e��hP�&`���G/{�KG�,�
���s�ѧ����e�r�7�~BIK���T��R���o�a�����
�FFVE>d;��)�*\>$�/�Z��T����NB��8�Gd�e��ŋ��tI��|�VO�X��u�v6�T���>����+�>����UC�	9�y��cd��H��f�

���reTO�@Z�Q:�و��Ȗ�'��ZqT՜�%~�~ݪ��޲���e�VX=�n��(8˅�'Ki���9�����
��=S��� ���XMפ�LX}1��+���6P�N�%Ќ�kR������pͬ0ݥ'۳����u���hx�A%��4�0�w������D���v�UN]m�t�>U	t�<dn�� ���b�;9z���S>�͞�=�2p	ɥ�n"?�_�@�F�ίHy6��R�-��u2�_f��������
��/D�#�Wp���v��,ѐ'��(�ŗ.g*t�o�Տ'���&�#�GԸ�@j96z�+'-K�r@�3s�������.g�zE��E��'U�PI?���&!�e��י�T����R%�W�z��$P��\�� �@7v��7�:,Q�VaN�@�*$�'p��+�ֺe���W��lm@ �e!D�%�wV�Ӆ�%F�S%��H�Pwq
4=���Xv!�0h6!��uL���[��yt4 �˻�V.�O��)]䌊m��M����hKA�>��ҚF�1P��23���d���:����3���2 �.�:,;-E0���N���E)�x�睙w&1�4�ͻ��{�l*0>��kMH�Z�Eq˨�J��4<~"�Va��D~�Ю��!��r�jq�Ϥi�aց��.�$�s�rC�B��&@�+��>��?Jio����d�
�KT"˪9��������.��(�,-��p� )���'y�����ƝRL2��%8���Ұ�a���8�c����c��~2�߲�0E5#2#?db����~T(H�1��L��9��Vs�/�mf4�>^
\�߇���+�vو�e���+u�;�jS�*$j�� ��*R���T��ĉ*wɻ�|d+hٽ�`hO��FF���@�d�/���!����`/��;�M)���