XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��;�(F��GE��s�,�p�	U�ԅ�s����~8������F�u*�
i�-��bL�Gh��O]��(�oo��$�ȃ�����o@���˺惭G�AJ�Äi���~o7�?K�[���qS�� w#x�T���/���<
h��~̱אe!�EJ撵6�S�)NAl����S|%�9V�iw��Y��<A�:������Qי�R�9�W�9ѱ��%x&��ׁ4
u�[W�t�F���y �쭡:!��Zb9,���X��EJ���],l�^�J$YiW��3L���?���@��-u���b�2�/�~�'�u,-�}ZjT��Oz ���J�\���05�XMk\�j/�-��s�C3���B݀4��-j��w��֊w�w�kȔ[<ux�����\��I�i�ϰ��A�����Q\S҈y�L3�s^�]=@�����H��"jk��8נ��Z"�vX��T	)����S�Oӣ���Oz��}F���&�)������4��э�a(�KR{�D���Q���^>�z�ø���o�*�-BĄ.����X� [���^&G)!�s�L���@������-��>�b!@��=���i]q��o�g�l��Q�;I)~i�v�JY��Z����v��qF��#�|�ۛ$,��԰�o��;�H�=�X>��&M@����f��������aE�K&�c�Z�w]�J�]�E�s����|ow�w;�ʱD���5�o#�"l��~+�0���XlxVHYEB    3a46    1050�:��e�o�":6f���x���#�� mk���!�I	��6�k��K��[�:�IP.lqv?]~���r���9��1K��*S.ºNfO�yCV���[Ko�,��ص�v� +�N�<@�!2L�~�y~�[˫�S��;D�0����kU�̿�y��B�y�qQ�{*��B�)�~����eX�K�ܴ�am��+�΃)��h̊��s�υm�2k������,~�H�_s�Oخ"r��+E���HG�sΖQ�B��~{;)"i)؊Ykgf�v�Ӳ�� =Zt�Hα�d��W՝|�=}a���'%}H�^-�tF�!4*��F�յ��b8,6���"�h�"o�?B� c�#�}C�@�ȡ��H?*0�B��9���w����I�!4�8:��8v���d����Y���Y���؃�gJ;�(0��J"D�H^~��g;%1������P0p��&�Ұ�yL�-[;LJ���
�3'7�/�ُg����i���&�i�/�j9��Q����%Az��b�p���Q[JY�z�e�>˂*�&��Fm�N��6E����p<U�v��ױ)~�	����̡$���n��U2�w��'����
�mpƾ�FT�?��C��/OzJ}����ە��`���2��Z�,ޣٿA�;u?�Kq�G�XTV8���fkr'}D��oUWBB߳��K(�YP��w�'W[~z�x�G'J	Q�A�n�<�)��K>)dZO��I?�!�-,M�mz?��|�W�@�`���T�@,�8��L/�����
e*<y�H�FF>����!���V�����|�Შ�XJ�
Q�r�,��I)�4����j-�#h��{ �\�l��m<[Ϥ��2�m�Sx톭P|vX��f�21��3�,��f�Z�N9ڲ���k��:O�YFyY�]21^�ΧF=!��?��	�,���	�bc���Dɗ���̓�j�dz��F�V�6@�Ap�r�im,S�����z|(�4'��5M'���AyO�;��4R|�2\~�	��b��p%������v�$��7��DmL��1�\�)G�u��w��fM��Z�����r����BW��4��6x��U�l;� Y꾛K�Df��7��zBC�%zk���T�kń�Ҵ���w����D��]-]V���!�/�x3oպl$�-z�60��&�h�����jKL��b0J&޶����H�`�衯kV�_�&]�1�%#u�����t�~kƏrŁ1����,#�0��g�8%k��"<Ô*^�����C���<������Hb$��_��49!r�}oE��A~ӟ�g�x���D�
�J.��pPoO1� IS���b������8X=�>�^ٱS���4��:8a
��lu�g�Z����j�u��h��.Ĭ<N�b�}`k������A�@sY�^�b��/>4�3+����ڎ���Nr(�1�/m�`��b�g��6E��X��r qFʛ/��`��z��$*�!�)ᕻF��B�I��E�\�Y�ey	�'/T*c
�J�v]v�R`�(�;v�`��0U$����|M�Nelb��O<�5hG��o�N�����,�q��1
�(�dc�PW�k;F�`����[���ڑa��
��}6,��ꪪ>*��>{�	�=�l����-0�
_�ɜg0��m������H(�/!!�T���Fk�>�m$���~��Q4Y��Qӝ��9�d|�RkuV��1�p5u�'sc�P0-�aB��2m\]�s	�(��Me�e����ᒋ���#n�e�+8�2}-E��Ј7�Y~����\��;�=�*.��[���w������ �1����ft���2*�͟�a�����!7v}5:���4�;]�f��=�jˀ7�\ߖ��ow�8i�Gyh=V�hL6u�Z�sQp0UMGA�W@�B`�]-�z��,�jlԿ�I��#<��q�ڶ���J`^���}�o�Ο��b��C
��MÃ9�bA3v�7cs�A$����! `��	O��Z�\���N���h� ��R�"�r�O�i���QRPI9�m�����N�CodΥ�X�iyy��"Ǫ@�w�Z���i�hD�|�ڴ�	{!%�[��3 Ý�]?��ML��*/�s�EL�r5��Y$
 �!2[H�w�����̯r[^��UݹA�HeT��*�>$�ԫ�:?Z'78=m�<B��`��OљbI��r��Y6=�c~��#�F݋8٥'es1AKbam��ֶq�DN)��AZ�rc���9?�L��-/�e���߃��0�*J	®ӛ�L<���(Y̕A���@6���&���u�|/P/�X�E�J�R�<�͂&��������M��7��l>������ݣ���[��3<��	}</�C�I�y�O�)Y@s���hv����B�v�=3������:UJ��*/9'x#ߌ������ޔU�P+<�֌�M�YJ�f��B��H���z���c���֞j`�~���7�p�����(ףR�#֔q����VA��mlzp!�}ҡ]ˀ����ʓ�	ɾ�m�ѺⲊ��5��1��&o1�M�PIFV�9�s1�lT4����(׭n�uB{x�9�|�M0m���/�g&��d�!�$�Pv%���!�������1� T,��2&ʷ7_�N�]�BFZ�o �ᮞ�2~2���`f�6oB9cS�5l���O�0yA8v�!h���r����3S��̑�?��쌳�ńa�@c���;/�~�������ک��.8�s�5y�M�E&��%]Ar�/��e�FA,}3ZΣ�r1�	� ��&AFڥ+V��[�|��y9�b2\�@7��|�։"+Y�ž��P�|����ٖ'8׋�rW�z�z-�`�4p�}hج8�X�y{�c��^��Z�R}0�6��DB���eN$�Nʎn�@{��2@o�醶��4^5VW^�`q�o
�	]I	��Wr
�u��"\n�`'���M�$�͙tYq_=�T�<�����2+����<6R���n�0�b�O)���*)l��t뽸�ET��ēg��`��59�k0M��X�Yc�?��CC�����1^.����" ь����d�������:�,�i�q�/�L55?҅�]�����<e 70�h�E�\�~s8_v"	��'��L���:>�X�,��".T-x����U{I���b�7#������~�c1i��G35+E��t�j��	���x�$��~Q��߶��&Tu�]�Y��W6�oĠU��4��Ui�^j�`���τ��
�3�]=3�-��;��ف ��������bԓ���-���p%� A	�7<2�G��tpe�;M6���68a�M�*��5�*��a�S��P�K�ʃa8���'9قo�L�� '���Jm�Y: �h������_�2�4@OA� B���]����E�V�-��:L��G��eveC�Nq�S�V'�j��ܹ��2:��]��*�}���l?j�M�|:�ƍ¬�<�Η���H�����f��{cA!(�;A=��V\J^K��l$WH���VՓ��7�dn���'a
>�a�tTH�Վ�r9fb&G���5�2�^-	��-�u\�ls<7�l?���b0�����pE�pʁ�Q-Ԫ��;u��\�(��H'@��9"e���7�_��\�QkB$ao����r�� #����C4�:�:lSS~�#<����&��0�5]:�b��P5:�Rɚd9�����'�k�[�wv>����<�:}]Qc]��3�!���D&�v�r�;�GU޶�	Қ;Km�=;��|h<������H��<�~�t��b��u$��/�̽ �n�����bh����rn���b��r�ݱ���T@��'�>��KQ�\Q1HM�5?K��:\@�Ta����|���E�?i�?;��o�T�t�0��Y4��a(��'�����h�1��0�C)O�ɬ#@�Bhf��4�1%QkbYCܴɛ�_���g$q�89��\u ^���g�<}F���٪�7�N�&��;����#����o��ѡ!�3ɳ���:*t��n{ؕT�xj�@m����tԇ�^���i(�	�$*