XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����l���:sJ"�Q�r�zڤ���lD�([���K9�Wpr~�o��m��W?0�B�ᠤ�~wh?lJ�L6dD��up�J�� �#��p����\��^�i2z�����*?�C ʢ���� �c=��5w��u�5!	~�4��]#>t�.6z?��aK�juz*�rI��#m�ڑs[gޘ����:d����T�Y��O��T��b������e�>�-7��Z@��\ )��4��_��g2�RXl �Z](�\�~9g�M����޾�E+�W�b5x��"�VVH�j�����ph����"�dbk�\�sLh{N����V܀�ۄ*/��&w�4r
�?W
Uv�^��`��3���l�T3ˆ��繃:���V���6`�o�.�΀��V���� �	�5��vlH�B����?���ފ^|�g�u��i�(�,mK��
�xh �i��G�%���+�{�π� ]�j��ݡ�C����K�M.E��fP!�bx5�T�U��|ڗ0��2��9ԊpV��B���9��tx�b�',f:��2b�|Orel��_�˹�,��=�1"�Ȫ�(j����(Lo� ��]D�a�{[�7���\깦��I�&f�q��vK�{�fsEdk��k��|#@ Ůs�h5v��.���x����V��_-|�J>�$߯i]8�MjN!B���d̈M�v�*��$Ȃ�����8
��bv���p�w��눧+;�C��X��kp��-�0�J&��A�����0cz�+T��+�D��q״�XlxVHYEB    3fdc    1160=Y�c�}0u�n�w:r�>�/���n�0P���LV��(�? ��8B(F��b(����^��IՕ�Nk���������+�{,��:҇ą�t�o*l[���:4�Ŭ�^d�|aYy,.w�(sp�����[�l���r'�r�+�,�j,�J<k,�]hL��iDC$�6���H��f5�����";S�L$Z͂ XA����+�-uFFO�M�s�֢��P�2P�Z��Z���V��d A&�k>��e��������p���?!���ɤ�1�׵,<��}΢����6�x= b����-1D�OL�b�W��l�b�c麰3�>z<��SQ&�t�c�H�"+&��q;Tx��uҟ^)��	�E?�n�����"vNj�A�u?�j��#G��R�w��u��&g5N�i#&�<CUI�6�RR�٬�٭䃍���'�
$4r����i��6���T�Ǳ='{�}����p�!x5���$�7�Pک�).��D�M�g^F*xP������~`�W>4mb����2H✖[��U�7��/�8h⌠�_@.�7��YZ�V��E��E��( 4^WYvN�����)~�*ؒ� ��FbcJq� ��+��3P	@/�#��>�dG�l����ӓ�᫕
9��A�3�v�,��8&[��G}NR#K�G
����\�ak���H�/��QԱ�X�L��Y�CVh��}#�c����B��kم2r,����	q@�I�����S�G�)�K1��;�M/f���:ԝqP<���-p��錷�L�ˋ��C�P*=d�_��-��37���i'���Z�9O�+[}p���%���?0���*Q\�X�PVC������z�_b'�3�b��B�+���pH�KVlT��ˇ��5)�k9@�&P*�D(�|�@��շ2c0 m�+�����JG{j�S�no[�%����^y,Tv�T`��S8_�06��ų )��>��������JGxW����׾(��o�� k���J�A��0��(����XH���ő��`�kUk��t��V.0R??D����D<�O-���_/C���ɖq�΁�
u������-��"�u��#d�^)�Q�i*�)�~��#��~@=�j�/T��u�|�Y�ӕ���7��5�8j�:fFtO8���H�k�^(�>K��P2�Q1�$�aj������1l��RKͤ!͢����U�.�
.���%�`)S�f���t{���=�/V;�E'j����7(+$�w2w޾�2T\ҝ��]30������qE��g7�#x���ZR,��.�!�%`8�S����|���f�~�/+��af*jѿ|���ŕq�G���]���ؗ�u��\�lB~�t͆Z:z��a��0�9�$J^�A��Z�7SB�V�/u��H�-l���ko��(���Lvg��ݺ�TO����C�dF�f������~D�h݇���ӝ`�,,�)���v�>ć�	�fB� �,}2�%�Ct8]�Fݚϯ`�3�t0&s*>
�T&����NcsD�g��s�%�o������9��$&i&帒�Z(���G�>���R���=dv�i*ϺI��\
�i�\T1uC�����n}s�o96��^{l'�EQxR�pm���4�	�ti�,�\3b����_27��u��U�����_*�����)�Wn�j:��w���z�5(��`r��X�_���#��I��G�*Z��<��;�;suT}��lQi�3n����������Ά)�e��j�v��Ћ�dŽX���'�'�+�9�G�HCqDt���N�Vm"�~�H9%"���aD�}9=�\/�(	׍{���|�D�������`!���F��emN�DZn\E��Ԏǔ\����*T�쎸��C���L��uɬ.���
�p��8"��#Z��c}��~�M]���CS0{V�ӳ���C%�)��7�S^��I��▬�<�k�,���Uª,����7U�2�?�&�6g�u����
:��Y��d��L���K�bĴz0��~�6}]��;?]pf��0�&�kcY��!L9ɟ�
4t�!3y�ړ���Ip�g�2`?`�s$UF���Np Wk�I���7�a��ކ����d�W��s��c)j�A췀�M�؎8��c��$���e�*EϠ������L�t`n���>m��7���V��l�ǎ��^��^�����}i��E�ͩ�r^�����6^�6�,��:?b�	�@���:	:3<�	8/�� IV^��/}n�o��(�=�W2��MC�4�{w0ڙ����~��4@�V�z��Y[���Ow�'��JV T�͌�k��W����ŕ5�/@��`�Z�A؊X"@���U�`�>d��^)��v7j���|P����Wgu�ХZ>CF̗dG=L��H�`6	R���P[� S�@�$'g-�]X���������__��7�;e�������G���ړ|�cG%d肦B���0��d�/�@'_���F�o���tdR�K0�2K�W����z.�ӍB�%�2��9* �n��!��;*s訮�Y,�5ܨ~���f�����?n:'#\���zDZ���+�e�|\)ʃ�
oa��9Ѹ�$��&f����H��q��օ�*7�o�J�+9|y���G
>���¿�=�~�"&d_�WܛX,qd#S��6������
��! �'����*��JI��*����J~�q�+��E���	����<�t#$=N��D���%��nrpb����2�m- ;�l�T����1�&�um�6yڥt��
P@<r���*�+�0�K�$�4�z^tz-'��L�p3.,���:�	�|8
҉[���n�I������	�g��)�}�?���|�g��[�X$}�Q�����Z�_&G��9�*N#� �t��	��L<�I$�:Y �C'{�������7:W�=�?;�D�\�~'��'�Q�xa(@EǇ�svL7H�D�I�t�	���	f�!������q�	u����o��Nφ�W�	_�+R+�G��q��܆c?�l]ࠅő�ϊ����J��{)��i�o��ԗL�s�z�����&ٞ���!s�����g?�(�����7���K��@_�6r�\3��T�^��>�&���z�V���N�\�����3�D�^f�w�y*��"�{�"5?�-���=�hE�B�3�4ڑ-��xt�����Iv��!֨���N����+?�7�����[r+Ь�����w����ػlM܏ix}��ĕ7���=۩^�� �����*~�)����(���/��>@�����x	�P�Y�D�*�����U!N���z��ҝ�2�S�\c��4��C��p��Ԛ���2�MR��D,��H��j~i`~
��!$	k�7��m����ZB_VE
��`t=m�P�?���)����ߨC�םE[[^�P�	|����Y�f����^������v+��h�*!��G@8�2d"�P�F�z�1
����_��9ґQ��z����.w�&�}Q�{���	��1�:�R��r�3w��-9�r����ZM���{;6��5��>%�p_��r��V�)At�gH�L ���+DM	Z�oԾ��Fdj���Ң�XԖRL�'��.����}9P#�ȉTU�Ɍ����ǧ�?B:rtve���
�|U��*���&��|,ŉ2-n���<�#]�D��/���kFu�n��Ln�3�>8J_��F�jj�L�W8RR<�A�B�Ve��D|�g�M?�W�8�W��� ش2{��K!���>�>N�D�d�z�T�P�M���������N9_X�1��gC�)��6�gƖy'�m��Cc��ܰ�*�(�w+�F7Ev��$$+�v�#F���*gĜ3Cڑ���ΒF;Tˎ��X�c�׍�*'| �-w�Y&W��$``�u�#2� ��M�fLt��N@Y��;���w`�M�*���*��oz�_J��,.�����6]G�?Y��tll�ѯɑ�i&��ۙ��l�[PT�@ql:��K)�5NA��umF6��Ly���_��:�^(,=T�'�8��!6��L�$/��񯈕�R �y`��Sh��v�)�6߄���5zr��H y�_r@J�3G��w��&;�}�9����;f�,�U�r�em�6ߺȧ�ɢ �ں�o?SF�7P����nO��U,W�y�s�:���!�'MVpow(��"L�gV�Mh�7�E���J#�ųU@�UY��j�M%:�iN3ы�[Qs*(p�\^,@�
�NCN�h���a�5�uA�PI2��s_Q�3�6��B��WN��^��lt�W�/�