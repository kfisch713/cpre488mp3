XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��dh��T��͎����`?�0Յmj��s��q1a��0]��q��9(�ڝ���9ʚE/).���2<��˸[,[���$4�b��:?��b�dpy��/РYBM-�s1�%��.+�Z�}�'��U���X�a����9; w֯��މ%`�'���G�+Ma���5�����͸}6P�����7Z����&�oY~t�+���E��A��/HB�"�6L��.`�>NBt|ؖ�E�m��m� @�JH�I깴�K�ne���ú�[X1�i
�`�EcW��
lũ��K�������bn$�~ �hWV�M�=��!� ��(��$2�Ξ���^���p|�ᆂ�@�0�%�����_������\����^׺\'A�_��g	�8�� �PHJ����5��l�S�X�Gy$z���I�`��4��!F�p����e�����<5l�����hap�\���[9�
2��Jiw�G���qn��f�C*��Y�L�j�3��Z��B�[�=��T`R`E�N����g+ud������K�U��L�Y/d�B�9��y���5I�W�&s�Bt����*�|���Љ�G4ۢu��|�Hn���[��CF
(�P�ZE��V�8-�䢢�f�uG����7,3+E�IV����x��?G�lFR6w?vo3@W��0�p1����Q��~W�D�`�Aˢm�����z���cf�A�
��NEc��m��D���	����6�s�=��9(����릥��� �ПXlxVHYEB    3d1e     fa0�������{H��������x����X���`�t'��U���/�SS�*n�nd E����o8.[E(����O���S�[L�'��a_1JC�`�D���̨w7C�ڀ�]��4��aD�g�L
��4iB����7��I��	�o�2�
��T��'7Vs�F�2����X����S��8@j��yiU��D�L7�7o66M�G�] v��RГ���P�Ow^=��s���
���I�n�ɧT�֪ ��E����S75����%�=�VBn�Ey�Q�]Z���%���}pV�>��1�!�j��q��C��vr'D�F�N�X��[\$�U�Y�
m'/4h[�3M����w�VKGfȻL�i�Le6v����k8TS!�K�o�+.<���p��������l�ʖ]�#x��#2JU��F����j<Qa�������{������Vos�iu"�����wU&�3�Ą[q�����}��5��G�L��ۧ�H����:P=�/�zWg((kYb�ܬ��*�j��o��(���C{�!�\Z �����y�.l����B pM{��v�b���(j}f�bh�R!<��(���>��88{P�u����p�Ŕʢki��;ŉ���#�]qxǹҦP����E�]f�o	k�S{/{���Å5�k�%���jPێ���K��)͛쥯��Y?��ߐ��9r뮷&6᧲� ~9����gR����!��~.}Y�
�Y��
3�����?0�b�a�P����5=?��^%Ù��Э��GW)�&�{X�8_����m~HN��e�u�X��M���5�-��*��t7�S"��>��<U�1N��v��9��!zÐ�Y�y�:9K(G��o3�>S*�x��כ(���-��7U���I�����ASG
R������1M���(�\�0�E�l%�s;��,�]GI�f �L���݈E�<� � 1?(~>?��:Ld���'M
u�m`k�,6�����m�d

d}�� �-v�Y������K�Oxd�Rf�2F?�L���*P�ڂ^����Z�V�L Gј�)%�P�ZJ�<ya�'9��v�@��SVź�5t�vr(�`��/h󿕒I=�+���ǥ��$]Z�`FYWbڐ!���*����y.���K��wyx0I�S�u4�A	��\:^�1�R���w�O�
�� ;��ť]��l𣷶{���	X0��yꊣ���캶� ��@�n,d+��}�2�v7�f�P pȕ�#ZRN��Iy��0�َe�4#�=�J��(���ض �xDw�;9bR`}���#�0�c��8F�*`�>/��cO����ט����J��͎�u�oخE��8��=m�Uq�#�ʙ�����/�0��;��x�D뢯�ߋ��5_}8hd�Y�}�ή�r��v9�T���IC'O|<$�!� }i���U,�tPX��[^ѵ�~!h�F�i��6��/�ڜ�k'�mߟ�X����iuف������i�}!�b!?L�h�K�ǰ$o�5�(��[ %E��Oc�O4��̳	�����������l��>̡L1�S�*��Nn�H�eFl�"J���U�)����K�����1)2;تG2�F��8�V�r�tp�\x�<����R\�2�5�X���Wj�_X��D�^5�VZ���Ev��۬�f؜$�C�P�*����ABGɰ��sĳ��i���m	��P�w���A�j�A�Uf?Q^��\3�H�)_Tƃ��(2��cBz������a�MJZ�:2iP}G�P��h+�
.;90 ��c"��G����I�^[]f� 	��w���`zϨ��w�P�T(�:�I�6#����ԁV���^�)��\�v���t�51�I��NW>���5��A��q#����!�i�#͘RYM]��j!t(W��Z^�U%R���X��	R(~H��&�	u�m��������x��5��]�f����yS_.8l+C20��A��t��>|��O
{������柳f�<o��8|�.{�� ;��f�vs�B�s][%)�5��Pl�y�_P`��y����r�َ�6�>n��x�c&Q%��U�6�D�ԑ��Vqu�ϸݱg��^xq�*�(,D�X���0��v�x�_1�5i`e�#��,�=D)��U�ja�n����Y�(�X*/ =�if$1Il���
�������"L8%a�m&��k�����Jç<�!��2X�b*�L����XՊ��,#��ό������uyL�gv���2�x�#��N�bV�i��v%U�%@�&^���/�D�2���zʵ�3�@�7a���au'� z�(�l��F!{��"$xI��)��f�
����L���Q�k�g2T\Q��	År$�e
�`��ĝ~�b�%r##k��dK�K�F��o��l]�AW~!ݸ_#�)�=�})����km\��>����Q�B��8~&����1EN�> �nE�0i��ë��k�g��u]�9��e2pk�����.?.�+�/d�nN�a�PC��9��l��_����i�����Lf�8���;��7B��J�Ī�r^���df�`���[(�ġv�̧6��1��]�w�v�D,�;��q�r��Qɺ"wEAj�HHz.�*�E&B����o˦���C>��<���
P�ɿ��g�XA��A��Aw�o�E� K?<����_�K�1�u%���8��°�J���d5��dA�Hz����;�|B�S�ګ�#f�J{je%M��)�h�dtUN�;���zL�]�[���*d���N�G<$-�ˤjv�����0U�W4
��5wke�B��g���I�=�!��n�0�VGy��v�]o�i��)˴�����s�Dn�1�/��sB�+����s_���Z["��'N�R�\�ڤ�
pҁ���ɽ�}-\U����i��r�J�O��C�9~�,i)��k?�$;/��p��:s��t�V��(����`f�n�"@@]�㍉	���z��>����>v��]��Cy`�r�ؚ�N�E�r;��D,�ª�	��%��g5W�v���ԫ��o&!��� ;��I��&�~����J
h��#ɼ�Qɴ���i��&�,Ҁ�H;8�1u�)�Yz2F�D��Y���T��NL�Y#ğ�T��%4�����Ϛ��D_e��\�!�1/-MGX���ɯ�w�G���H���F�2�uLr��\��-Vko�����b�-�	��;��_���Ǿ�K���f���ĖQ�uˆ+���7*�3��r���t�����VyAז�/�����=���5���=�Q*�^H�
	��G�+�t�F�GqPQ�H��d�&ޑ�Z&ȥ�iX�y�[�^�K�I�o׮!\�Ԫj�����$�f����h�}Lji�v��`T3��N��~��ʷ�*u'�l��.�T�:�r��8p<��c����m(�N4!���Q`wu�`O����9 kٗ�q�S�gHx�P��b_��h���{=�a����]�ݐ���л �$�n}2����s��ݰj ���滱�"L�:�0�$�i���p�t�(fA9~�9�2F>h��A?(+����t�гڠkF�����İ��N4�T\��$q*D�}8�f/�Vu�l�5_��˵�͖�D��L��e��QQ" 9�I;��⛘�sO�mq��D�x�����'�+_K0�o�����=c���A��O �a^��a��Pҙ�q�!�ŭ�Ym��lJX�C��8�'<��]����fG���׀�4� ��{�m��b?��(-[�Ȥa;�/�,u��^*C�,��� ��� ���WU���-`��U���@u1�<
@O �/���@������mnw+c�id{Jt衐�&Eq3_���N�@tUI���}W��0X�v�q/H�?��