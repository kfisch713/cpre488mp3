XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��D �,2E?(���� @�{�������0����������߯��/���=���)��-�P\�d�����+��+�dT�/������ӡ�:����H9�apCu��f"B��2</�B��gZ��[�b�Fs��J% �*?)^��H5sk5��^\_S��jCi-n�(c�:��/JR��:^Rf��Jh�L�ұ#�n�L1��d㙺���h�y0$],1�`py=�L�G� �&q�Ğ<�ΦV�D�6��n"��:f6���$��� ״F&���1�&:=���o���@
�ȝ�����t����;���ꆱQuL�?�`>�0�&e�e�kɅ{�!6U�����{8���:P�����(�HE����?b|]���j/#(���@ϧ�L|��s��N�(s��K/I�<�0�ѱ�����q%6��ʩP<�{��6o=�l�����׿����YJAm�>43�Q{+iO�W�R]���m��n����e	Ү����'HL�ƪ���SX�f7vF���iY�PaÂ��7��K�￢YB"�й�ė��&��7ާ����6�Ջ� �H�(��yL�S~s��HY�W����#K��Q���1PM&�n���;�
�di$�m���^$#�>�"��q 1�n;�����74s�OX	Y3�4T;R��|�K�g�v�vS�>tO���X�X^M�b"�7�u7+je�E*v�j]Ϯ���+��W��DnNŖ��Ѻ�{3g���S�,�=�22+(�ŋ%XlxVHYEB    3a46    1050�{�r�]���~31��T��[��${���ď�EFl���ܬq��A#H~C�� /�A�m�(���rЁą���P����/,�h�|+`�X|�TT^��u���{�*E��7����N�����u(�zZ~��:!����P
ϻ4��="�'Y�����d�v	�,q)S<�� �+4��Hm'4�nPi�����s�u3}���m�f�!�}ѳ����>
bXA���n04����}���e�W�;�\��bu�+��L
�~�dܡC��{�*f�B�'�٥�H�a��O��:�
����`o5�|�pőYiJ$�ѹ�|�w[U.i������W�}��M�]S��/^)�C� �2:���a~��_�$Uz��\ѣ�e]�*���7�&Lyϫ|��r�R<�_��rrX��h������pmf�#�d� zq}�Vx��_�s��� x]N����]��N���Ŭ�+��V8|����'h8dp�3b���N�%`��zAG�%�_u(�� �Y�j�g��QhQs��|���Ꝉ�?�QX��}��z�nV��'`:d��!�E���^�8�ow��A9ғHُQ�����PgJ�f�)<��ײ�5r��|�芳�
��A5!
�3�+�֘�R+݃��ښ����[=I��A�$.�ڋAX+_��j�,u�)�Tn�w�����Ra?��Ͱ]ܪy��b�(ɹ�8�>�wh$��O�Q#�r���8�u�mF�����{m�����!��s��HEv�O��5�V���W��>��[k�1��4i�x��B�����[��)�f�[���o�8�?k��m����Ltي����l$��P���{�{ъ�?�Ǚ�b\j�i�<@���s(VR�K�@.��kmz��m]
����n��e��Bo���9o��
�-:����[Ҿ^Z�Ԏ4��Qh��V�[���4*���6ˈ�fm�\�P�
��碣d���w�ߗ�٠��{峹�lC�3�($q�&f�K��G���-�.�����*�0��l�����\�Bv	EN]ڏ 
�
�(_���^���RH�ٚ�n��������#�1�+�Wh�#���C��: I*��;�|'�"�tD�N.,e��򈧈6�1%���+�wv��ڿ�r�|���I�����֫�Z��][��Β��RH~���<�D�L�{O?�[:>���fP��e#��N��� ������\yb��M��;N�g����G���S]>H����ozȐ��6����] t6��FA���˃L��Z��2����i9"�!\/��L�F���mq��彟��h�`_5"�	��s"X���Y��[5�Dmm��ٸǘP��ÿNم����P����ez3|]Z����U�t%)�&�iY�6M�)W2*Y�	v�	ں��_��'v�&)S����m��4z���i�v���\��cN�J����l	Cq��xɠ�eJ1F�gC!3D���BF0P�I�+B_lY�R���ux7ă�~���������+/B�]8��)���������B�=O�jV�P�?9�O�I 1�|@�d��/��:R(z�j�49�j(R�������}��?������׫����QwcB�SBR0�Fɲ4�K���j������	ˌ��=�}B��P ���G?�,�-�o?����C�p+
��.���p��O͡&�#HY�>+�3A��! PFc�v�/��ݍe��Iϥ}�V��3��)2�2M�I%\�X�7+$pHƭ[*�|0f�+9}MC���a��3J�a�Q-�ֳϑ�ʫ�XC�Y]���;_L�o�]&�����M�&����H-�����x����]i���4v&��&֨�E�/�V�)[/�~*���Wg�����$��j���*�H.�!Z��ׁ���k�":w�u}�Y�Q��F�RH�l�v���b&~�&tʀ���o���G�L-- &�c���-y�f{�U� �٘@x��j3UX�L��<m�i���YC推j�i���tw��QA����X��_0��6�?�5�g���������Z�3n��-��8�R��Vޅ�Tg͚!Sk�G��޷!���Y��{�tm�+]�H|Y��y"*=�������f
�m�l���Ûb/)� h~^�����pNV��>|�ψ(	2&��}��Z�@Ҫ����{��>-΂����=4Ӣ�ǻێ��G�� #���]ߝ�7Q�@LV�S�I1h,N��'�U�x��m��z_uV8,bL?w��d�D�~���+\h�h��ص)��%�];d^D��Ϯ��z9XȄh�EK0�]0�a�;����My�K�p���P��\���#&�3ӿ\�x>l:��А����a���B��Mv׆e�������5�>��`A�ޫDTЇ�<R�Pw�+�FO׶P���ەŶ�����CаH9j��Te����a@��[�J���a�́�K�r��i
�_��cF��z��n��ۿ;�ǔs�1X�}�-$���ipf�./Ö��"63G|�[d��@�'��U��"ʛ$�ge�'�ѵ������L��Â��ɧP3�w6N�ɻ�sR����)	�#��&�W_��Yc��e�Y|p��[ݼR2g^��?I��2���Z�V	���k4�3���Q�Y���=�!šbb��<���ky��Mg�f���2M��>M$��K�.�����8�Pp,���zzc!�!?|:V.w��&��UlXl8lF���8�~�y.�_7�_�P1C5��6�d�z?LG!�ȿ% \!�`9�y��Q��֠_���"	�]"��.��Z �SFg��!A�i�Xm�%��5�	G�����E�
-/!`I �1��٪>j"���L��-[r�y ����� �����d��8N#}�;.>���]�?-(�d�Sg���X��'aO�9<M����b��]�}�,���IJ��2��@���u3B���K���ZJ�J��O�-���e6B�$�Dt�9�������L����>=��ߴA����q�n��j�m���z�>���s�B�S��7po���`-�hD�p�o8�\�*8|ﰂQ��>�5��Z�y�'� $eyl���Z�,P@R+)�2/|$��Rb/�L��C7�
��g6p��#k��0���7���~���m���D>?�!�D�6�.CtO�:��]Cv¹�U쫓�/4@:�W/s0lTY~9���l��3��V2�k�)w��2�4� ��2�/�fq������	��џ�BQ�?�FuD2+��/˪�=Y���.���c���{F`�-�hWZ�p��y�A�i��f��qa�����i7y��T�R�9!�C�4`�=��� �*�AӭX�������0�
�J�ɽEh�Q�h)�//�cP~Z�:�K��6;����R���s��a��l��;k�N��(��8��L��Q�W�ޒ���L"kM�uMpTpW��Q�Cq�_pG�d�T_����!	3P��Y�̖�d�U"3��}�I���G���
����ρ�t8_
�$���	!O`ؘ<?)��PeC��ukO��Zz�������D��]�[*���*�Y�c9�*��P]̅-c)���2I��� ����sɭ����;��rX!�^�8�/+$�ER����&�E�R����y׆��plڤ�y�˽�(�7�3shO��S����+�\���~*�q	O��[�P����`0��#�LY���Ԭ/{����і��Jֹg��)g��,�:��g<XN��x{��o`�2�
H�ȸ��ր�Y�K@C�j�����b����&(�|]7�����G-��x�ۖ�_0�.�n*Fګ������*���'I�Y$9����diN'[��?2*3l���t9�(�2�I��+�ܤ�2���2qli�I#ЪP4�6����6���f��}a���:�ӄ�k�p����0\~	����yv���_35C,+#��M�s�c�߉(�V�h�e����
�귯3`/�^����
&�P���>랹�+z�w��4
�VG-�Nh�*7-�^E�*�Z���77!S��:�ə�~���my5�缳ʲ�'��>q�TP)�v�m�$l