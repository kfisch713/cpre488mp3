XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd����t���7ad���8�������0`Y����e?9c��jm�Gdk�1a	��utffO����o\�sV��px�=TG�zK@�ׁR�aN�zg�9`��h�
��<�$�(�P�6��E�S�nU�Us�V'}'���4��_�S�)Fye#�0AڨH���c�a�~�*�Ϩ{��W4>3Y �m*��֯]�liz��\������^�{���.u�
22��p)hft��˘c�j��S�y�L�FS��7�ׯc�\!�5��V�Ur���yʨ��ƿ[镘�AߙIڽJz���Di�1�'�t�J�{��ݚ@8A�����@$���qq�qQ��.564L;R��M١�7.�]�:Qkk�1+�ƀ��lj �g�Zݮ_ l�5�S
��~�
l��������b����9������"�\�j��ǳ��[Nm���R�Z�E ����s'� �	@�r�g��7�(/t�D�͆�p��� ��-%��Q��u7�t~��+;�Χm�e�T�4G���3���'�8N3���gsg�V�D����ۅcF��J��2�{��/����)�JӋg��`ѥ�j����tn�����#��E�;dX-�w��<I&W��vq&A+���T������+s�'�F,�%�N�7�<������u�7K�:!�W�GG���D?��v�qk�������V���-���
��ǌ�h:|��ZNf�R�3�8�����q���/�R�8�IW˩D���CXlxVHYEB    5866    1100���*���X�"YE��e����>�� 8����������@�[^<���� wi�7��b�<sM>�"t��iR�_�ȁ8"�Ve�^����B1W�=����D�T������6�h�T���I�D��_�0G?$�L��+���C7(WŘ�+��[��^����sd��I�|��X�}&Ui�&����	_I�?�6�BZ;�����u�s'NX�?��^�P+ X�Q�� s���=�6�乣��pM�3I��ɰ��52�.w���9��~/�#u�����.�G�P� ���#*���qc�0�?��[�(q�z�xVm����� ��06r�K�:�����P��$��e�ϐZ��e�U\~6�/�$��q �<��>C�A�c���\+�o1���+�M���qYg�Ӻ��]�^�)�ς�;���k���d�u��u(�ECk����D2*�w�xa��N�l9*HJ����*t�?o����%x��9X����ʳ�yǮ�塚K\���1Nc�wh{*i���`y�������h�4��P��(I�Y�X��PqvMKH�*���v�d�}4��x�o( ��T��=yގ����А@�Ռ����s�����y��<C��.�殙�;0$R�T�C����S��Tzt����ՍH����0�P��$&.�3*�2��}�rb��}9����y>#�*�=vp��[1Tz���Z�Ϫb|O�>)etg��S(��Ѭ8�����76������I�}L���c�Ne����*���vl����(�W�/о�v�hֵP���M��X��gA'D̩�TX�O�d��-��x�xY�x�~;L��)�M���ϣ�2��d���C�>�|W+����j�a��LWO���l�5?��8�ݥ�AD����k���O ����R�N�ڪ��g}���$ۻ��>��"�B��58O��C��&/�EU���m>��T�ώ��H�s��8�l[��:"Y*��C�d��#�t>A�e������p�g�Y�����Bغ��[��B`6M!N�n,�Qxj��Kչ�5�"��8T��p�����;�?��wLn�E�+�p�%lQ�n��ߩ��)�1�z�u��b����OH���6(�I,�[8�ʦ������RlC^hSB�=���6Wy]��Q&p4�����
���\ʹ���UV��t�/�m��ğ�U|k��|%>�I��ΖR����w<��$�en���G�](�p�m1����Mk:f�G�}��7@���L��M��wE�g�7Ð~�3_����sv�PG� �Oף��;np���Q B7����9�'���S�V��������4,o�;��`�_�>�h���3�J|՚��if��8d� n��aW2ױ����t�j���o��^��Ą��T�8���~[�SB�Ll޲|�>���^����pdF�B���PzW�}�?�+	CG�.gc��9cTJ�|g��?����ďngG/_���Ⱥ9I�vn����3}�6��[-��ne<0۞���ITW8��K���q�r��f2�70ݖ#�P(��Q��=��CM��>0>⹚��#5W��Y��M��"�X�`Y��9(7���=��t��ŃF&3�f��[��X\
��/6hYgN��;l��˫�{�������#hA������P��_�-�S̄ъ�`:]��}�CaחW[���S� �ş&VEŸ��>��`�N����O�={��ʷ0;�#Z��g5��f�4g���R�@�p����"Z��a�9�r��_7s�X����B��.�r�+V�L-%O���0� Y#6:��N$MB'7�0�(�t��5+��bN?�t9�w=���)�,���ž�|��;������-�}$T����jl� \!�Z�����|�v�0�H+k(b Ex�I̤� �z�n�u�A�q��9������#���(�$+�N����)x����X�����8�-r�$���ɴ�$�����y�\��Pa5?`f煆�����V��F�;F����98q������\���qt5���x���H��X\��wX��"(��:�Z֨4����Tq:������x�~�Q�t�8�.�S����%���`���M�
DE��v�J��t��O�}��q�r�穋����(�'���>��<�e-��o�誎v�u��C��ÍI2�����MH��$��B>�(�˝-�#�LF?(�78�c4!�@����١��zͻQ�۬~c�JG�tIC��<Ho��{w����=������D��zXm�i�0����:��ً���@��?Xɩ@�n���p9�����o�Fm�'_D������PR�(�q\T-�������j��e��	10��,I��������� 	'h��2��G��f-a(��{F�X�[2�$�'��XLPUf�`7�^F]���/������+������ i����i�����JNEȱ�����N��}'FW�n6���Hh'��Z9@D��By�#:�:{�a�j�m���r�����/�0��,f��6�]���"�S��{���ͫ
��JY���uPs��1 3}��������U�Ko[����Y�{��������s^E��/��.�R$'�h����:yt�������|~z���߿g1���ޠ���b�f����5��Ύפ�k��L��)uK<\� ���a#fқ Fr1��vl�N���՘C���CE�M��LMl�|$��ŉ�((rn��l�ȍ���*(gj��D�����bG&���s��0�-z~�K���x7c��J�f����܄�Գ�k���Մ.n9�J\L�X�5C�N/B�ۘH@����eVG# y��lE� ˜�ǵ�\BϙO�r&����4���6\�Qu1Z�9��j*��h�نRf8}�-
u�Y��X���M��2��T �z�I�1�s�G�Ǉ�/�<ѝ��x�k��g�-IB��'�:��=��@�o56�d�:$�;����9�I���<���2#iK�4%:�5�I�������gY�)ޞ͹�@� 5F����W�mh�,7A�f�˄�C��-r��3�H��x��UG�D{O�s��$��GїN��"��Aт��CQ!���$����7��8)
��U6�g�Y���.Vc3�qԙ}섚�i0��D�Y��H�Xz�w(���;{�!T٦3ʽ6p��#��v�b~�n��Uk��Vu=��J�ͷ�>m��el��o�I�<�ϩu5`q�%�A�U8�	7��ry���"�F�\��.� ��D��Ro����
��S���s��35_�e����~�yd�|��.�/�#aF�R��gІoG��Z�Z%�p����2[��J�c��w���6%H�rA�^���ͩ�x|�)��tF�n\Kp�t��=bU;��&���/�$��'_�"�Ϻ��>�h`;M��.�l�-������)ҍE=L�Gr��~}�i�a��8�Ttޒ}��=˃�����\A�i���FZN�%b�|ş��1���@A���J(���¡����:�f�0i�!K���7�ۅ$�Dr��*S`�ؿ-��	H"Id������`~�Q�mq`�д�k:L;0���gp�oc_Zh��Zh����t�
ܦ�]�H�z�������T@<��N:��pָh��"���K$Raڕ��ꮼ+'[�W�xKYX�!6�Ac/�Ey��a7ED3�;��]݇(��"��߳}��I����od�f�d�]R�t�����+?l�s���m��V���- ��I�sl)�5M듻D�-V'˨��Jm|g7�����l���3✇6&����*5��>R�
�c��l`��M�J��hH-ܑ��!��돑�-FQ'M�AEl4�n(����tB�H���r�ڳ���;<RNm��Za���
�R�����tE���"-¨�	 ����q{��uk�H���졄n`��?Y�{�D��Nђ��a�����q�=���X��,�\UQ�����G���u����t��t���}�0M�r{՘��e��vZ��=v�i��V���5g�� �,g}gB�j��2�}�>�����!��z�ss����6�n�Q:������F.�����f�����xC��$-��9�lWpC`y�H�f�8�m������+L�w�0���5dm����v�	I�o���M߹��1��q!�$ 9�hp���rt����!RBOF��6C�|�w