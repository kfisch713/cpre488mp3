XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��AP�pg�\���*IY%SN���m�u2��|[��ؤ�9Y Sn-�o������5�S��vW���O2� ����(���2���>�$��]��v�"܏H�)%\���v��X�8۷��P��;�/�_L���E��
�`�'�z���	���Sk|`c�"m�`���H�=L�� +�'yp�|�9��+��I�T�� .����}%��[JC��u�{�%��4|�T\��y���$z`�l�v��S{V�4��y���[&1� �mȞ�����VN�5����ES�u2=^t�Jŕ�d���(���-�yP��P�WxS��B[�1UAb�5A<���Uџ��I-z%�(��Π�H��wB������5g�ϓ�Q��U^��乆*�_pޱ,���57]�8�v���$���?%��{�*��-�FU5�\B��b�A�������U"�̊���M�unM[*#l������j���x�*s�����e���5<t��%.
4GR�g�'>#�0�Z�
T������YWy:�υ��+篪��ڋ(��]{� 4�BW��ВdA/8�=��Z�&<�Z��8� �`��y'@*{U��a�|mq'#R�cO�.�E�a({~~f���������+�X��M�To���KK�l�G�}7�8�׆���=u僝K�#����b�'Ȣ�4c� M�	��O[!}O��i	}��K+#J&'�)3pgl�{��psڊB��e(��	��d�^�i�P��NFq'Z�.a���XlxVHYEB    290e     af0j?6#DlA�V����~0�c�E«}���F�iwL�:��?�Do��ڝ�����T���n�{샀1���2���}	^�i,��T�a��x����
���|�ue���x'Fp��漯)W-̜zxG�0V�S�}N�ƫW6���9�< ����&���oW?@elv����3�*黏���,v���+��ġ
����u�{��G��Z�aTzH���"K�#�I0�÷ug��Wׄ��	�������>#�
&L�P�k'�@�����~N��0}f}L(�e�r/d�h''L[��L��b�I,��c��5Q�:�B���L��v\њ��b3}���S�5)��W�o'.'	҄i����� _xE�a��O���*��+��2�n��C]ܩ~�������_j�Gw���i8�m����O`����V��8�ҷȘ�Kti�$}q� ���zp�N���q"�L��^�c�������{|����6⡥�Ħ*�orl~<I�0u�l����^P}ŷ�T;SV=�R�4։=D4�D,]�U�,�@�۷���0�Mt3����^�˵�8Y�"��PH#�luZ6�e����qg� �v-�^N�.�U�I����>�:=�;�H��i��<��;`�	���T��C����
@���"3+�۔��k�����V���p%rDO�B���
�kw3{\,���b� 0��G��� �����n~�Y;�K�9��w��X��e=HQ6+zlɛ\�l~��Ԃ8F9C[��>rҙ�P�^�G��U�'W$��gB�UD�a�?fS�]<c�6�y#�"lSue#�E�eS�I�i��1��a-����Į�ߛ�rX&.����� dY�\b�7{3��,��|L؎�0�,�2IK�mRO�(n�9�(�^�K< ���=D��yiT�I��Y��_!�QyF���k�e~����}�M�uۂ%9i][d��$��k�o��ð�,��iN�=�点G1�������ڽ�c���ň�0��u�����F���)��$R.�X댶J�#���U�:m	���[>��ڤ/��p 	\3�o�B�(r.� �������� ��&=��J�$a����~v���dm3YSc�G����;�����| \�;+���po�?�"H%�н�5%���{������X.�~����S�$Ɇ,GN/N���L�G�XO�~�q�bN�6�;y��/9����	�q�W��;����fL/��Z�"nC�F�����k��XA�O�D��:^���?�餣s�.���.`eEN���n#��\��X'(�2�f�^�eZ�tleH�W���JJ*K��9��-� ��"O���#�q����*�����"<��R������v�/�=bsR������#�M������w�����o쳭Y��9v�1�*���Zg�Ti�9���t��K�3����d�5ٻ��h��z��k�����3�>�V:����ϯ�3��X�w7���LȪ.7�T��A��Yn� ��土���`T��;����h�p�
��m���wM#9����<�@���S�8b&O�RR���~w�P$ c�?� ���O8��jW��@��g�n�K䰐�dq�:�;G��b����!(ܐpV���%9>�@� Z��v
 gR�O��D����cjχ̻�s�M��u}����I�7@�>�0�h ��
Q�O���SHF}�Z6C<��D���u���)&f��;/jT�~
�%��g\��ܣ�6�Ɵ,��6zTK
h��H����dc<���X����T��3MOZ2B����ES�m��4�?�∨����J�U~P��ȋ�]�4s/�c���byD�����h�ƒZ��\��u��%���e�k�l*��${P�Zm`,�,<'ʷ���.Ԃ+p�_e�s������6��t`�R��э�/��*c"�xz���$9T.�922������;�tX��J��ʿ�֊;�_*���KT��i]��=��J4��ҋ]nsRk���{!��������p�@]�(���UY���>FFGV��-�~$=u�5�xl���.yB�_�D[���L���]� �jo��f��HkL�ռ,٘?�Y��$l' a�,˄8f}s�&�BÂ3��۪�sϲ�?U�05s�Ro�`VMB%��s!!���}������o*f���Ǒt#Q-Iτ$I-Q��0�N��ܹ��]�z�a;�HD�������:��a"̯�!$g^����hpY��%���j�,�So��ӱ=�������ٵ�<�m��h�w "�20�DK���b���~r��dL���!?��ؚ��3���{ɯA���y�:D�Y+���m�Y�YWG��ĭ<5�G�:q���q˩l���c��{<�w����^��jL �g�N�''F�c�y��	*�2}c0����:���M�c��	;��k��U>��C�^�t�0"����p2rK�N�b�%#�ն1��^ǵ�ҢuQ����	x���_ e1���v��z��g�|�����2�8&aql�t���.�7԰&��Le����&�)���B�%1.V%��(sa�n|��?xsg&��G�y��ى�7{w�UX�L�
V�����z�dΏ�
ݷ���L㵸.?o�����"<����2}K��		o|�lX���3����O/�~M�Š��i���@`�_�l�p��P,U��O�t_�4<�I�`X6ヾ2��^����[��N��a�Y��X��fV$z