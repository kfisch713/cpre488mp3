XlxVHYEB       0     58c��$+w,� ~3�8�ЋF��9C�s�2��0x��Z�7�[R�ht�:�a�b�y�����}b+������������]�M����U�������D�:YT�Eϐ�'�m����e����bO=�M5X�E�DzA{�M��+���"�F�9��"W�k(S�f�w��&��d�#,e%�N'��5˴�H��,�G�e��`�Q��է|�x7�ue���nb�ưy�Z��~��'&��Nہ �������OȘ�Z��+n��M�{a���Yt:7P�j�y7u�������Z��gM"�����-�Q(/�(3V#�
��HU��y)�x�����Q�_�\	�
$/Q�-�͓���[��
z4�D�	���a�����ţ=R�5�D�Bѱ��8�<��v���f�h
N�wC�ʅi�D;����#�to�W�{�l����-|h���㙣,r �|��dx�=5P�3! lFv�����-�rF���EJ����_}��M�`t�)�CT����d����N��ß,,ˬ�i0��Gk���%�X��ߪ��;�PI	�!�C�$r}�Q03rI��2�VP���Q������
1;����'�KKgp��o��q�yd��Z](�Q��Z� ��#kЧ���,`&���a`+Cv
��8T7��JmY�]G��
س��k/�4�= V7t�{d˩ 4Q����J��q�����@�QuHYi*Å�|��sn~�@(<|	��&��l���t��`����	��Ĳ�������`;�.aZ"�w6�a`a@`�b�jg�w6aMf��ي���~ORΎ�����H4,j�Ae���,��%����(�oo�[�&a�vUovW>bz�Kv�q\�+N_�8Ir��G��v�X��^ wb��0]#��h��'O9�D�fѺ������	��Χ_~��E��$�T�Odb3H�3��@��9�^8&X>TW��O���d�.aP�?s�@��yr����B��F��~���B�je|E����i2C�\@7�YC�U��jO��?f�M�6)�Pͬ��c"�¡��2B��A$���\���F7n�d�l��#��i��C��X8���`�R/6aUӂ�̣�Be��{92��6��ZuU�W����@h�0֋�O^I�uV�����)�м�:���&Q���z=�$���6��Y"80_.�MKJ�#%� ���)𪹷 x����$Z �R��h�h����5qg��uM}��l/�q�bA�U�*Qѐ#8E�&r[r���'����'¼���^d�-�)�8�6����ׁ'�.9�p�����`�;
����TqA��S����;ܱ#Z�s6���e9�� ��bY����ok ��(���e�l��Ӑ�H�P�!�XlxVHYEB    1421     7a0ؙ������S?�]ZJkJ���⍈̓���X��j{T6�Oz?t�e���+ܯ 3u����[6N/�����	�/��������j`u{�ݦ�i�,Y�'@�Ǿ�ٽ����}�$�f"���N����,���
�M��3	�O7ǹ8 -Y�<6n�0? ���V�ʍ�2���"\b�y��ׯ�HI~xv�hk�v%�#cՓ����`��1i����6RZ���Q �)��Dj�vn�h�kٚ�w�K}�벅N|����1q����Y���T�k0��2�*��pL?���"n��q��.��$�Ĺ��Ͳ��M�q"H�`�<�^��&XlD�IY	�ࣥ�Xh�	���/�'�&x�	{BfZM1�@�	�T��<�0���DG���r`�����dٓ6?CgM��'�䗔>�b��q$����;Ƨ��������[5#��� $�p䨖�t��*V�:2tL������nI~�S���<S m!B��}�>�8N�\�e2����t���ˇ��d^foK��ѧA���S��XiB�h���l$�Q�w�z;zo�y�xR�[H���C�	@������i��+�/:|�#r�X~0 �5�)JM�%b��e�S�@��!q!�
���.�*��?�Wbt���h_��;=X�j$����|Zx�((�S`�wKY�xDW9r ���ө+�����ڸ���Wu�K�Э-ؓ�p~�%s�qs��!� �.�Y
��T�6�̴VX�rn恕��<�6>���V��ߖ �.���o[�!�����0�[���{bT�
=�l:j�c�h��jnMD�th�RL7 ��u��s ��J��B�����%1���[���0�����r� ���)��G�5�-,|	¼R�i|� q��ʆл�1���J�;�R�u�
)�����m5��{�-�{:���N�Ԡ�P�GoCNQq	���g�$���35+Ц=�����";!�
��V�)R��˞�f*^���NL�z"B�U�&Fw�vZ2]2V��?��F��v���f���"�g��g�J�Lyb�w���e\���:Z�����3nWP!�m*$���Նb�`%����K�;�!�]G���&�+8L%]�R�lBD���rZJ ��U�,s����7{�'����f[���$��x�6b�+F�y�2��|
d�4�|l�����C�����s��I׮��
xbJ�����);w8�]�D�f���(#��D�ȼt�j}#�K��ט�/�-e�����Co�Tґw��u1B��gZ<��|�v$�v�!�#S=�6I����y���j�P)�S����n��\v{̬���Ԫ�B7S�y�	�����Z��xg���<zxв�e���b1#��?�����f5kF>�:��]��tEl(�Lx5�y��j"椀B (�X�dk4�JI����L�Zg"-�~�?%��V�f�,T��(Ǯ��ĳ:�%���x=�Aï6�	]�=>�[2�-)��	��ap�5�L���3N��N�wU-�娺T�U�����6������-
ʶؖN�~;1���������i`#��hF�N�8��������"q�H�`�8^�Ħ�p�i�|�6{Ba_�_�٨�0�oG�+��H1�����`�;:W���Rdڴ+'��Q��_�;.C�;��]�$^��~x֣ĺ�O��0���C r��?��9~,@"�K6-��a��$��v�`=��4�h�T�C7Y��#؇���$a���Dz5<t�h�p������]DE�|���&�*mcLq���tM��_M*�?^��J��P1���a(��z9�vwn�X��cG)2�p=�܎=��j��p�Y��YN�O�!�c⒇;o�!��L��80l^���6��44�; ЇҀ1s�jY�.eƮ